`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bditVpm7Pw935qRXUQ1sETq1+PglaLBd+aSPYeW88FSoUtCjxQWy5va7mz6h7LJIziUYwBwD+j3t
+VMSP+slf5LjUhxFAKLks6InMEDLndfD7RWTu+fOhUvdB1FifhbPzW+c9L0tAH9vCLVfrFLPq7vl
yf4zwX7oVA7lqmqBAP6vjviH/oy0uJxBRrWbc5tnB6MIhk/YRmVJbsJ8XTWGk8AjB/GYBqoL+wpq
pBHqjhuplvzds1RUGVbQcWCEYb84XQ8jHW/hF1U8BUx9miuwurgqmCmOQ3xJmUjd2rows6Y4ohvD
HnuNcWkjk6imR7+MFucwyQFnFKJcRW8RZBcgpA==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
S9D6gb9IpXUjtHQ2a6AkmOem4UNKagoQdDpwl/Bm9bJF7Gg0+D7N/YX2KzYmBCbVj/++hH/MXjXt
2hb3eHLoSQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
km3Afrr1suGsyNc1U6UnNdNRISFGKFeFZbegynH2sAJyFyFy9o9kdmh7U7D01FlNDpoK6sRCVTa4
eJBk0yr5ndP8iWQprTjeVsl6/Z0TWQQ3e1BgI1OJE+nidvJEafrKdyLVunWOjG9BZmqBpRuhbDqm
bOFBGPEKeaOrO3NjPSY=

`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AbEzylMLdX46giKSnq27MCQdv+o+LuV0+ZeIRc/oFQq6vAli5csauAGMb3IS4gHnnnXZyL7YEZYm
XHrh5bBe0SVW+RyOKoDK1XMkskgptLTm1bGb8M0rMZRCwxAPEIs8y17bu5Ge0FBFC+9ZEtvU/zEn
M99SqmiM3V7R0L6qHvw=

`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
G5LuirAbPHZrFevioFcRVQFYB+49SSTOCXKG6dabN4bai+MM9/ZaMBASMD6DtCj/t5VB4NqFRAYs
gTHPIcd2s4wmfHOuIymuHHYe9aV+RxPwAe+yRU5wvca7QO8trbsGsUlgIEsm+uAt876MUW6SlHrw
UEn7G4QFYiibTOUEWVYMimVSZSEmQtLtxmM19qzsrwFZU7L7qI5UoNS8zpFPPulaUT6ueLJHWwDo
blVV/tdB4cT8YIhi+Mrw40tRo6Uz4cZMzloN3WT3CKGMlfWTXwJhWzO4gY20hx4UNbT8vIAfCWgj
YzYT0ub4v3FX7TvXvc00Yijtw9Sy9NAXIt2dNg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3072)
`pragma protect data_block
A349HNwWYkD+rVoCssNnMONs3v0K+4XVnlsZEqu8AFPZxl5u58jEOVo4QezAuGupeEoYu613N5Ru
IBlr1Qf9MRJD4CShzr++YOeNwB+opYFW5F63aWfZWZPFWqXRTAPRszLcvKzD0Sc9LCpuVP2NSqfa
tsiStd6u4r/divTTNuR0HWgmDcQMnlUsFyaVpPJxhbAT8tpeAZsG4eB0uYfrGirJUwmneuY88dkj
CHO9c9goSRGl+33vKJ8jQS1gHpI6SfEACBYbzpOh+nOD3qfAFVvIuuV3jB4Gv7/BYkWcJmxbLYvE
s7VTEIUVGVQp9sS5D+idfukYXzXgiiMed3sXMp1rJgQB5xmaW3pFZXrRBCzYM0jfVN1nWfACga06
z8UXxT+9mydwJuPIeFtVKBPPSUfSZpJPvC4i5+2PvMZPYRnVaSJ/ZkbYZR9Oa8Dg0SrmIsYCLCU8
xoFZp9W1SzHYM2oxjwYFpRZxvzAeOAzoBn4/Hy84Fg10BtIG7ZkXzONNH+jevCla4UVIP9cUoNY5
8Lg0qzyOXZMEXRU5KcorGmyNcON+AULYpi0GwYuX9fOY4QVp3Q633QddWSF66CPvBhQTU54RW1L2
TcIAIdVsJ1v2Xwm805xN58/keq1hHJ2ZUdc+SvqDyBGiylE6599JCqyCJY1CrfdskTUvw0DBioST
89MOI4z6uXfB9RVwtmGE50M8FuCKrvk16Zj32pD4wGlwb1nqwA4w0GhV1hxWgxqaKOB2R8DtM3TP
/LymVfMxxKfhU4wz4sdTUDdK3ozZAm3Tphvqub+/VmecVLemBqfJtPAJjqPnwc7TTc9BoVeubzSr
UTWYDjEK/l9aVLpf6dyR6E87AYdp/u/3N/c0yx1Cg14FWbv+oVa/gQbcZpdVIAUGgM8ILIxz76mJ
ZIkAKfq6R62O5Sb1eImAlLxBGpnyDCD/UpssIXoNPGcS4lKEP9zrWZf9E1xAZW/MPu62qMSkokBi
Sf2XOH2+xap1BuEJfzn6Gqq57WXOOCcMT7fs+4C9PS+o/QdF0wTMdFh+XmoFMrzBrVvCYbneu6JP
WoYBUkkKippSJApX0hNYM0waS/gaUZ5qwkiiC7eDRukQXMBZKHw3eFRhp2uvAf8ab9qbujuYgGr1
w84IEZCa0oTEA3G5EDPLWPZRRYbqNqB2HXnQLXFVYl2FQR8GzkbA9a665C7kQEZBZyQXDWGhTVDM
H//lH9s7X4cLCnuPjgeDJQpNC8b0lbDwWzHjaEk/dquvGM0ippTKaFUJlE7vv0b+vvi7UXjJkWIr
wqBzoI+S/S/NuQO0X1PnWkoo3DtH6kFdXGiDDfZUMM0/SoqlV41lij1vrxHlMZY2hpPoc1VBHGBl
pjfU9DnwGjHtjLFQIjC3ByIZN8oJR/OZMnxj/d/nNPmVoTmiIims1saLKhN6mV2ohin9xEBNdtem
8eSi+BcicpprKboNq4HkHfOPkgb5o/42Jq5fEf19ZQAn8iOg7Ovxg3OaWA4vFXqeaHBdNNV5dDf2
295VmlkaG8Ob9qRQhOgPDE6jLHAUoP3J3O5gmRLFD93fTCmVYNap4mQDs85taqpMyBfJh58hlvB3
1VrOWpGKTXevBjTKqWQFW/RZqz9+/EXrN1GthtfGSalwmm8B+PjkdwRPw/Du+NSP0fmu/LVewPa/
6DBzguzuta5GXgdRG1tvfrUsWOsDrazoJNb12d/WGX0lguEz5ybXZJNvYmnG9ApElMUZKXab8xnp
65r8edjwHEvOE8GLeVkyfjq15npXZkBKIqALGJJ+MXzLozZ2VFnrzTzcCCe5NzmpGLmovrSBuxo9
7n+7EKgDgR5xuKqzvdCxj0BLxjpoZm8Fe+Hcc24/cWqq889zhMT9Z9xZTPgx5h5rLRs8x74Ye3ql
XBykCgZ1/ilsxVF2sg+0yWQfww6oCeZdrFuixyvRkqd+ueKMMpv3fgsKjOqHjJ6WSiEsoCPYHAT/
T6SFZ3Fj2Snb+eBRe6Jw/+tAvnpHT/kxo+y1q+pxg4wVf76GyqGuZjUn4yhjIiOKv4JKhTd3jGer
JoE5siiXwDnOKTBr6+3fcZ9AC0qz8W+2dYAlR1bUjxF/vRIO9zLZq9t3fs5bJnQvFtFPx5CekVRi
9DgpcRhWcibldOX3OF1HTQabtQ0p2X8VbJSgmgEJNNNs9rIjPFt2Z8e0mTvw5axlgzPKlATVT3Fz
7rNxJwRiB7vl3VeC6SDgiAlCsdZ6TsjiAf9kRcDBhKyy68p0W982C5yUfSELibzf7DjKG8UeIxoB
N4eZLd1RAtcPaYa7C+ej4E2y615a5bj0iJYklSLvy8ZzCPJrtCvn/X2djTxIXONiq/wvh1DXc7o2
UDLHaUz5NfG0x7ddxDPqS0NDfYt4uXMarBpN4720f20fQqEaMqJM6NaQ2rnyLX7xnussqQhg7/zE
TKd8FHENFNYgZXuXUanfPSk2gZUOnuFO0iO0V23ye1JtvjZ9r4ZRJXaWpmRBX/G8YQ3I7LO3l2cK
mr3j1GowkorSC0Z1lAYIICH9Rmk1JlHVKqslJ3UlL4oYGsBlFh2VRkXUAMAdk+Qb9pdOouqs9USA
/TWDaO1sEMEV14sslTipeedUGmjK5WcDyRBm8tYzLgVkom009s1Zt+3aq4eWyNh0q7wy5eA2ctqh
JW1U+On2N06c76cGH5Jw234AxF+Lpn20WMraTK0WvuvJe+JPDvMrj3GCt9Zx9tnQXvyYgCaV+QJ5
IAmeq0EsRggks8q5oQHxNCTyhjnAq4+UgWTfzSWfFQBQe+749KOjEJ0ChtMPUVX5jieWn7VFoIPF
x6ykRty08HtNMWtZGYVkTLlvo5N6i5oZ9k+LqnVpRrCnCveHpZLsTLGVPS1vOwTaryki9yKEQ6vp
NAWQm6nJcbRHyPQ/UHDx4sA5lacf3ZnqpIR6/YxSATUkDvcOYCfU2SP2h9ccj+4PpomB2s4Xb/g9
bUMa4tEbuC2fbD+a/Z5BCksYiiGOP+taYjPiVoZ48XCIIZ8cNxqbFydxUGTBlzJuQAd7AT0v7r/D
uqXTwcTbwm6zu3hbHyQkFKq0PZa6gGrV3XiLvBbOT/yiticILn1i35bwbRPadPs5ul9GupjKAtw9
Egdu/WnBdlBuVyQTrRWozdMiUg+ABVEPHGLHN+ulA6kDuO3reY2upbr5SVgygwKlsk5nCcOnPfXP
ZEy/ju0/93mDDnfI1dibVSiNF8BwirNyq0nxle+rHL/Mnwd6u7cZqCuxh9Ma3642/+ZmaZhb+n0W
GYCDcIjvJX6blZAylNCN5H/DY6aljCg1XDWak1IAbTJ6NGcASwHLlplFXgCGTDYAEn90Og8V976L
CUy3dbBs+oIMbYaZwSwHUqH0eDhl+47G88jq5L/Efx5yg3WqEOqCntKqv8jixHAySW0OVX3FEqq4
z7s57YKhMmi52MmAb1uetUemTaspyJTXaFehRhwZpY1wE0rlJ4/kI/yOPsGwiyRKcYebPcmgxLf1
V+Zox0yQ02fN5iDG0aI/sKSOoiPmsUf3ePyD8AxJoTFY87Aazc236hmVn/j/ieYsIK8L4o/F2sau
PrTooT9wWRMClG/024b9yqnUSpVso6WQNns8rRSmVVFZhzkHHDIzESZPxtntzcz0vUFkqYyGcFD0
TUiwKLrl/NaKDQIrYyx8rANSpApbWS6MsKPggrD2DokFJd6Cuj6fA2D3j+Ik3QASIicgkcgot6b2
f4MAHiGPOFQgT3D+a7I5zSSdgs15OPOLM4lfJI3dKSutZHyAEBzMjQTzugvJJ/edNDbpGQt8w6df
cj/myJBo5WvUpwIMa7rvPfZxPjdCtzTG1O5bAz6/nxNvIbqdvnW5da5ofJSjSq8USmL1fIBcThUb
6g8FYq4aXLT7OUX/cwthjsfxbDpmoSFyan7JZDbR6yhmtz8ueV5X76/UYSIzOu+A1uDFe5yO1r9f
QG+5lKGY+84EAbgb3IVAhPDkESfciLbiFGSPkJAyN+A+8fpBy2zeyYyKE6+yKi9UqE9VrErgBLkp
MT95znS2EDGr65WOTKeEYHLnKDC7EBq9oSOUBjN5IdvpU7nGznwcsN1D4La+zOQKO/46
`pragma protect end_protected

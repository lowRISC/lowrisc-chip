
module picorv32_axi__pi1_opt(
    input logic clk,
    input logic resetn,
    output logic trap,
    input wire [31:0] io_reset_vector,
    output logic mem_axi_awvalid,
    input logic mem_axi_awready,
    output logic[31:0] mem_axi_awaddr,
    output logic[2:0] mem_axi_awprot,
    output logic mem_axi_wvalid,
    input logic mem_axi_wready,
    output logic[31:0] mem_axi_wdata,
    output logic[3:0] mem_axi_wstrb,
    input logic mem_axi_bvalid,
    output logic mem_axi_bready,
    output logic mem_axi_arvalid,
    input logic mem_axi_arready,
    output logic[31:0] mem_axi_araddr,
    output logic[2:0] mem_axi_arprot,
    input logic mem_axi_rvalid,
    output logic mem_axi_rready,
    input logic[31:0] mem_axi_rdata,
    output logic pcpi_valid,
    output logic[31:0] pcpi_insn,
    output logic[31:0] pcpi_rs1,
    output logic[31:0] pcpi_rs2,
    input logic pcpi_wr,
    input logic[31:0] pcpi_rd,
    input logic pcpi_wait,
    input logic pcpi_ready,
    input logic[31:0] irq,
    output logic[31:0] eoi,
    output logic[31:0] dbg_reg_x0,
    output logic[31:0] dbg_reg_x1,
    output logic[31:0] dbg_reg_x2,
    output logic[31:0] dbg_reg_x3,
    output logic[31:0] dbg_reg_x4,
    output logic[31:0] dbg_reg_x5,
    output logic[31:0] dbg_reg_x6,
    output logic[31:0] dbg_reg_x7,
    output logic[31:0] dbg_reg_x8,
    output logic[31:0] dbg_reg_x9,
    output logic[31:0] dbg_reg_x10,
    output logic[31:0] dbg_reg_x11,
    output logic[31:0] dbg_reg_x12,
    output logic[31:0] dbg_reg_x13,
    output logic[31:0] dbg_reg_x14,
    output logic[31:0] dbg_reg_x15,
    output logic[31:0] dbg_reg_x16,
    output logic[31:0] dbg_reg_x17,
    output logic[31:0] dbg_reg_x18,
    output logic[31:0] dbg_reg_x19,
    output logic[31:0] dbg_reg_x20,
    output logic[31:0] dbg_reg_x21,
    output logic[31:0] dbg_reg_x22,
    output logic[31:0] dbg_reg_x23,
    output logic[31:0] dbg_reg_x24,
    output logic[31:0] dbg_reg_x25,
    output logic[31:0] dbg_reg_x26,
    output logic[31:0] dbg_reg_x27,
    output logic[31:0] dbg_reg_x28,
    output logic[31:0] dbg_reg_x29,
    output logic[31:0] dbg_reg_x30,
    output logic[31:0] dbg_reg_x31,
    output logic [31:0] dbg_insn_opcode,
    output logic [31:0] dbg_insn_addr,
    output logic dbg_mem_valid,
    output logic dbg_mem_instr,
    output logic dbg_mem_ready,
    output logic [31:0] dbg_mem_addr,
    output logic [31:0] dbg_mem_wdata,
    output logic [3:0] dbg_mem_wstrb,
    output logic [31:0] dbg_mem_rdata,
    output logic [63:0] dbg_ascii_instr,
    output logic [31:0] dbg_insn_imm,
    output logic [4:0] dbg_insn_rs1,
    output logic [4:0] dbg_insn_rs2,
    output logic [4:0] dbg_insn_rd,
    output logic [31:0] dbg_rs1val,
    output logic [31:0] dbg_rs2val,
    output logic dbg_rs1val_valid,
    output logic dbg_rs2val_valid,
    output logic dbg_next,
    output logic dbg_valid_insn,
    output logic [127:0] dbg_ascii_state,
    output logic trace_valid,
    output logic[35:0] trace_data);
    logic mem_valid;
    logic [31:0] mem_addr;
    logic [31:0] mem_wdata;
    logic [3:0] mem_wstrb;
    logic mem_instr;
    logic mem_ready;
    logic [31:0] mem_rdata;

    picorv32_axi_adapter_opt axi_adapter( 
    .clk(clk),
    .resetn(resetn),
    .mem_axi_awvalid(mem_axi_awvalid),
    .mem_axi_awready(mem_axi_awready),
    .mem_axi_awaddr(mem_axi_awaddr),
    .mem_axi_awprot(mem_axi_awprot),
    .mem_axi_wvalid(mem_axi_wvalid),
    .mem_axi_wready(mem_axi_wready),
    .mem_axi_wdata(mem_axi_wdata),
    .mem_axi_wstrb(mem_axi_wstrb),
    .mem_axi_bvalid(mem_axi_bvalid),
    .mem_axi_bready(mem_axi_bready),
    .mem_axi_arvalid(mem_axi_arvalid),
    .mem_axi_arready(mem_axi_arready),
    .mem_axi_araddr(mem_axi_araddr),
    .mem_axi_arprot(mem_axi_arprot),
    .mem_axi_rvalid(mem_axi_rvalid),
    .mem_axi_rready(mem_axi_rready),
    .mem_axi_rdata(mem_axi_rdata),
    .mem_valid(mem_valid),
    .mem_instr(mem_instr),
    .mem_ready(mem_ready),
    .mem_addr(mem_addr),
    .mem_wdata(mem_wdata),
    .mem_wstrb(mem_wstrb),
    .mem_rdata(mem_rdata)
    );

    picorv32__pi2_opt picorv32_core( 
    .clk(clk),
    .resetn(resetn),
    .io_reset_vector,
    .trap(trap),
    .mem_valid(mem_valid),
    .mem_addr(mem_addr),
    .mem_wdata(mem_wdata),
    .mem_wstrb(mem_wstrb),
    .mem_instr(mem_instr),
    .mem_ready(mem_ready),
    .mem_rdata(mem_rdata),
    .pcpi_valid(pcpi_valid),
    .pcpi_insn(pcpi_insn),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_wr(pcpi_wr),
    .pcpi_rd(pcpi_rd),
    .pcpi_wait(pcpi_wait),
    .pcpi_ready(pcpi_ready),
    .irq(irq),
    .eoi(eoi),
    .dbg_reg_x0(dbg_reg_x0),
    .dbg_reg_x1(dbg_reg_x1),
    .dbg_reg_x2(dbg_reg_x2),
    .dbg_reg_x3(dbg_reg_x3),
    .dbg_reg_x4(dbg_reg_x4),
    .dbg_reg_x5(dbg_reg_x5),
    .dbg_reg_x6(dbg_reg_x6),
    .dbg_reg_x7(dbg_reg_x7),
    .dbg_reg_x8(dbg_reg_x8),
    .dbg_reg_x9(dbg_reg_x9),
    .dbg_reg_x10(dbg_reg_x10),
    .dbg_reg_x11(dbg_reg_x11),
    .dbg_reg_x12(dbg_reg_x12),
    .dbg_reg_x13(dbg_reg_x13),
    .dbg_reg_x14(dbg_reg_x14),
    .dbg_reg_x15(dbg_reg_x15),
    .dbg_reg_x16(dbg_reg_x16),
    .dbg_reg_x17(dbg_reg_x17),
    .dbg_reg_x18(dbg_reg_x18),
    .dbg_reg_x19(dbg_reg_x19),
    .dbg_reg_x20(dbg_reg_x20),
    .dbg_reg_x21(dbg_reg_x21),
    .dbg_reg_x22(dbg_reg_x22),
    .dbg_reg_x23(dbg_reg_x23),
    .dbg_reg_x24(dbg_reg_x24),
    .dbg_reg_x25(dbg_reg_x25),
    .dbg_reg_x26(dbg_reg_x26),
    .dbg_reg_x27(dbg_reg_x27),
    .dbg_reg_x28(dbg_reg_x28),
    .dbg_reg_x29(dbg_reg_x29),
    .dbg_reg_x30(dbg_reg_x30),
    .dbg_reg_x31(dbg_reg_x31),
    .dbg_insn_opcode(dbg_insn_opcode),
    .dbg_insn_addr(dbg_insn_addr),
    .dbg_mem_valid(dbg_mem_valid),
    .dbg_mem_instr(dbg_mem_instr),
    .dbg_mem_ready(dbg_mem_ready),
    .dbg_mem_addr(dbg_mem_addr),
    .dbg_mem_wdata(dbg_mem_wdata),
    .dbg_mem_wstrb(dbg_mem_wstrb),
    .dbg_mem_rdata(dbg_mem_rdata),
    .dbg_ascii_instr(dbg_ascii_instr),
    .dbg_insn_imm(dbg_insn_imm),
    .dbg_insn_rs1(dbg_insn_rs1),
    .dbg_insn_rs2(dbg_insn_rs2),
    .dbg_insn_rd(dbg_insn_rd),
    .dbg_rs1val(dbg_rs1val),
    .dbg_rs2val(dbg_rs2val),
    .dbg_rs1val_valid(dbg_rs1val_valid),
    .dbg_rs2val_valid(dbg_rs2val_valid),
    .dbg_next(dbg_next),
    .dbg_valid_insn(dbg_valid_insn),
    .dbg_ascii_state(dbg_ascii_state),
    .trace_valid(trace_valid),
    .trace_data(trace_data),
    .mem_la_read(),
    .mem_la_write(),
    .mem_la_addr(),
    .mem_la_wdata(),
    .mem_la_wstrb()
    );
    endmodule

module palette_mem(clka, clkb, dina, dinb, addra, addrb, wea, web, douta, doutb, ena, enb);

   input wire clka, clkb;
   input [31:0] dina;
   input [31:0] dinb;
   input [8:0] addra;
   input [8:0] addrb;
   input        wea;
   input        web;
   input        ena, enb;
   output [31:0]      douta;
   output [31:0]      doutb;

RAMB16_S36_S36 #(
.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h28287E28147E1414000000000028281410001010101010100000000000000000),
.INIT_09(256'h0000000000402020364854543C282810242A1A1428585424785414183050543C),
.INIT_0A(256'h001010107C101010001054383854100010080808080808100408080808080804),
.INIT_0B(256'h40202010100808042000000000000000000000007C0000004020200000000000),
.INIT_0C(256'h38440404180444387C4020100844443838101010101030103844444444444438),
.INIT_0D(256'h101010101008487C3844444478404838384404047840407C0C083C4828281808),
.INIT_0E(256'h101000000010000010000000001000003824043C444444383844444438444438),
.INIT_0F(256'h1000101008444438100804020408102000007C00007C00000408102010080402),
.INIT_10(256'h384440404040443C782424243824247866243C28281810103C405C54544C4438),
.INIT_11(256'h1824444E4040241C702020283828247C7C2420283828247C7824242424242478),
.INIT_12(256'h7624282830282476704808080808083E7C1010101010107C662424243C242466),
.INIT_13(256'h384444444444443874242C2C3434246E545454546C6C6C6C7E22202020202070),
.INIT_14(256'h784404083040443C76242428382424780C384C74444444387020202038242478),
.INIT_15(256'h282828283854545410101828282424661824242424242466381010101010547C),
.INIT_16(256'h1C1010101010101C7C2420101008487C381010101028286C6C2828101028286C),
.INIT_17(256'h7E00000000000000000000000044281038080808080808380408080810102020),
.INIT_18(256'h1C2020241C00000038242424382020601E241C24180000000000000000000810),
.INIT_19(256'h1C223C2018241E003C1010103C10100E1C203C24180000001E2424241C04040C),
.INIT_1A(256'h762438282E202060700808080800180038101010300000107624242438202060),
.INIT_1B(256'h1824242418000000762424247800000054545454780000007C10101010101070),
.INIT_1C(256'h3C0418203C000000702020306C0000000E041C24241C00007020382424780000),
.INIT_1D(256'h282838545400000010182824760000001E2424246C0000000C10101038101000),
.INIT_1E(256'h0C0808081008080C3C1010083C00000060101828247600006C2810286C000000),
.INIT_1F(256'h000000000000000000000000000C522030101010081010300808080808080808),
.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
)		 
     RAMB16_S36_S36_inst
       (
        .CLKA   ( clka                     ),     // Port A Clock
        .DOA    ( douta                    ),     // Port A 1-bit Data Output
        .DOPA   (                          ),
        .ADDRA  ( addra                    ),     // Port A 14-bit Address Input
        .DIA    ( dina                     ),     // Port A 1-bit Data Input
        .DIPA   ( 4'b0                     ),
        .ENA    ( ena                      ),     // Port A RAM Enable Input
        .SSRA   ( 1'b0                     ),     // Port A Synchronous Set/Reset Input
        .WEA    ( wea                      ),     // Port A Write Enable Input
        .CLKB   ( clkb                     ),     // Port B Clock
        .DOB    ( doutb                    ),     // Port B 1-bit Data Output
        .DOPB   (                          ),
        .ADDRB  ( addrb                    ),     // Port B 14-bit Address Input
        .DIB    ( dinb                     ),     // Port B 1-bit Data Input
        .DIPB   ( 4'b0                     ),
        .ENB    ( enb                      ),     // Port B RAM Enable Input
        .SSRB   ( 1'b0                     ),     // Port B Synchronous Set/Reset Input
        .WEB    ( web                      )      // Port B Write Enable Input
        );
   
endmodule // palette_mem


/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'hfe0e9ee3fffe8e9300a00e9313249a63, /*    1 */
128'h0962829300008297ff01011b40010137, /*    2 */
128'h000005170bc2829300008297000280e7, /*    3 */
128'hbe4303130000a317000280e715450513, /*    4 */
128'h006514630020031300555513000300e7, /*    5 */
128'hff81011301b111130110011b4940906f, /*    6 */
128'h00000597000280e714c5051300000517, /*    7 */
128'h000046b7fd9606130000f617f8458593, /*    8 */
128'h240e8e9b000f4eb7011696933ff6869b, /*    9 */
128'hfe0e9ae30085b703fffe8e930005b703, /*   10 */
128'h0085b70300e6b0230005b7030006b703, /*   11 */
128'h0185b70300e6b8230105b70300e6b423, /*   12 */
128'hfcc5cce3020686930205859300e6bc23, /*   13 */
128'h40b787b300d787b30107879300000797, /*   14 */
128'h0000f597305790730907879300000797, /*   15 */
128'h0005b0237a0606130000f61700458593, /*   16 */
128'h020585930005bc230005b8230005b423, /*   17 */
128'h00100913020004b746d090effec5c6e3, /*   18 */
128'h4009091b02000937004484930124a023, /*   19 */
128'h008979133440297310500073ff24c6e3, /*   20 */
128'h00291913f1402973020004b7fe090ae3, /*   21 */
128'hfe091ee30004a9030009202300990933, /*   22 */
128'hff24c6e34009091b0200093700448493, /*   23 */
128'hffdff06f1050007334102373342022f3, /*   24 */
128'h6e61697241206d6f7266206f6c6c6548, /*   25 */
128'h61207469617720657361656c50202165, /*   26 */
128'h6f6c6552000a2e2e2e746e656d6f6d20, /*   27 */
128'h656d20524444206f7420676e69746163, /*   28 */
128'h636f6c65722070696b53000a79726f6d, /*   29 */
128'h6d656d20524444206f7420676e697461, /*   30 */
128'h0000000000000000000000000a79726f, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'hca8686930000f697b7edfda007138302, /*   35 */
128'h87930000f7976294e20707130000f717, /*   36 */
128'h87b30280069302d787bb878d8f99e167, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ea17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c927837e4a0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405264080ef498165224b20, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a2852222a080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000e9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc8e498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d924051c4080ef652240e050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h888505130000e517864a608ced01842a, /*   60 */
128'h740270a28522186080ef65223d0050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c398050ef860505130000e517, /*   64 */
128'h543514c080ef85e505130000e51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h120080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000f7977139bfdd4501808261056442, /*   74 */
128'h04130000f417f426f822639ca3478793, /*   75 */
128'h043b840d8c05b9e484930000f497ba64, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043379ea0a130000da1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h294050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c5016a1060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h051301610593460978f060ef00f11b23, /*  102 */
128'h00041323082c462147c1781060ef0044, /*  103 */
128'h00f404a347c576d060efec3e00840513, /*  104 */
128'h757060ef00c4051300041523006c4611, /*  105 */
128'h0144069374b060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398938787930000f797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h697060efe436f4064619051984b2842a, /*  117 */
128'h162347a168b060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'hd51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a0017ab040ef4a2505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef5a2505130000d51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d7230, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d0023551060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934d50, /*  146 */
128'h378505130000d5174bf060ef953e4611, /*  147 */
128'h978a350a879365b040efde0254e25a52, /*  148 */
128'h445060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a30320079346d060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h0793449060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h427060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h06131020079340d060ef47310d230001, /*  158 */
128'h07933a7060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13df060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d0023331060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb1323060ef, /*  173 */
128'h307060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232cf060ef9d228562, /*  178 */
128'h0000d51700fa2023478512079a63000a, /*  179 */
128'h0e8801090593461145d040ef18c50513, /*  180 */
128'hcb840513978a3504879364852a3060ef, /*  181 */
128'h3531470328b060ef014905934611953e, /*  182 */
128'h0000d517350145833511460335214683, /*  183 */
128'h00a146833501578341d040ef15c50513, /*  184 */
128'h352157835cf71e230000e71700914603, /*  185 */
128'h0000e71715c505130000d51700814583, /*  186 */
128'h01b147033e9040ef00b147035cf71323, /*  187 */
128'h0000d517018145830191460301a14683, /*  188 */
128'h01214683013147033cd040ef15c50513, /*  189 */
128'h160505130000d5170101458301114603, /*  190 */
128'h05130000d51755c2010157833b1040ef, /*  191 */
128'he7170121578356f713230000e71716e5, /*  192 */
128'hf6bb02f5d63b03c0079354f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a35048793371040ef, /*  195 */
128'h35048793359040ef148505130000d517, /*  196 */
128'h140505130000d51795be978af0040593, /*  197 */
128'h40ef14a505130000d517b501341040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd3330, /*  199 */
128'hd517317040ef13e505130000d51700fa, /*  200 */
128'h35078793678530b040ef142505130000, /*  201 */
128'h148505130000d51795be978ad0040593, /*  202 */
128'hb35d2e7040ef14e505130000d517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85162505130000d517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2bf040efca02, /*  206 */
128'he7970a7060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439c302787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930c9060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0a50, /*  213 */
128'h0fc0079308b060ef000107a315410223, /*  214 */
128'h025060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e105d060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'hd51785aa808261257aa27a4279e26906, /*  223 */
128'h34238101011319b0406f052505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h101867857ba060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'hd597842a000546030015468300254703, /*  235 */
128'h40effa2505130000d517fa2585930000, /*  236 */
128'hd597860ac10d842adedff0ef85220d30, /*  237 */
128'h40effaa505130000d517f82585930000, /*  238 */
128'h0000d51780826151641260b285220b30, /*  239 */
128'h095040ef1e07ae230000e797fc450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'hc80a8a930000ea974401ff05049389ae, /*  243 */
128'h0000dc1706000b93f98b0b130000db17, /*  244 */
128'hfff58d1bf94c8c930000dc97fa4c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h015040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057f6040ef856602fbe2630ff7f793, /*  250 */
128'h7e4040efadc505130000e517ffb912e3, /*  251 */
128'hb7c57d6040ef8562a0317de040ef8556, /*  252 */
128'h40eff22505130000d5170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d637c20, /*  254 */
128'h855aff2dcce32d857ac040ef8556a029, /*  255 */
128'h00f45b630009079bff0479137a0040ef, /*  256 */
128'h04852405788040efa80505130000e517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e90905768040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd75e040ef8562, /*  260 */
128'h86930000d697893289ae84b6f022f406, /*  261 */
128'h00009717e9c686930000d697c5096ee6, /*  262 */
128'h854a85a6e94606130000d6173fc70713, /*  263 */
128'h85bb00955d6300098f63842a6e0040ef, /*  264 */
128'h40ef954ae7c606130000d61786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c296c20, /*  266 */
128'h27a060efe4c585930000d59700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h0000d517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee6ac040efe3450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'hee8707130000e7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'hd51785aa690264a260e2644202091663, /*  276 */
128'h879346816480406f6105dda505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b2d84505130000d517f86102f4, /*  283 */
128'h40efd7a505130000d51785a2c8015e20, /*  284 */
128'hd517690264a285ca862660e264425d20, /*  285 */
128'hd51785aa5b80406f6105d6a505130000, /*  286 */
128'h481958d94781862eb78dd3a505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c21101df6808130000e8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h6105d1a505130000d51785aa690264a2, /*  291 */
128'h0000d51785aafb079de327855600406f, /*  292 */
128'hfff7c79300e797b357fdb7f5d0450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h8932cb2505130000d517058514590087, /*  296 */
128'hca8505130000d51785a2c801510040ef, /*  297 */
128'h64a2690285a6864a60e26442500040ef, /*  298 */
128'h71514e60406f6105cb0505130000d517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'hc58b0b130000db1703810a93020a5a13, /*  305 */
128'hbd8c0c1300009c17bc0b8b930000db97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h444040efc14505130000d51785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000d51785d6963e011c0ac5ed63, /*  314 */
128'h043b66a23e8040effa060c23e436bce5, /*  315 */
128'h557dd1350f4070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a23ac040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae327056722120070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h89aa04000613fd4e7115bfd58f8d2505, /*  329 */
128'hf556f952e1cae5a6e9a2ed8600884581, /*  330 */
128'h577d67869982e16ae566e962ed5ef15a, /*  331 */
128'h55796318a24707130000e7178ff98361, /*  332 */
128'h0000db174a8503800a13440106e79d63, /*  333 */
128'h80000c37adcb8b930000db97aa4b0b13, /*  334 */
128'h07815783ab4d0d130000dd1708000cb7, /*  335 */
128'h06137786028a05bba091656600f46463, /*  336 */
128'h77c20957926347a299829dbd00280380, /*  337 */
128'h04090863792227a040ef855a85a2cfbd, /*  338 */
128'h0000d51785a60397e863018487b37482, /*  339 */
128'h64ae644e60ee557525c040efa5450513, /*  340 */
128'h6caa6c4a6bea7b0a7aaa7a4a79ea690e, /*  341 */
128'h40ef856a86ca85a666428082612d6d0a, /*  342 */
128'h77a274c2998285260009061b45c22320, /*  343 */
128'h855e85ca993e86268c9d79020097ff63, /*  344 */
128'h2405006060ef854a45818626210040ef, /*  345 */
128'he7178082400005378082057e4505bfb1, /*  346 */
128'h869300756513157d631cb7a707130000, /*  347 */
128'h057e450597aa20000537e30895360017, /*  348 */
128'h862a0ce507638207871367858082953e, /*  349 */
128'ha00505130000d5178087871308a74463, /*  350 */
128'h0000d5178006079b04c7496306e60b63, /*  351 */
128'h0000d51787f787936785c3ad9dc50513, /*  352 */
128'h11417c07879b77fd04c7c963a5c50513, /*  353 */
128'h05130000e517a4e585930000d5979e3d, /*  354 */
128'h05130000e51760a2148040efe406ade5, /*  355 */
128'h05130000d5178107871380820141ace5, /*  356 */
128'h05130000d5178187879300e60a639ae5, /*  357 */
128'h0000d517830787138082faf612e39ae5, /*  358 */
128'h8287879300c74963fee609e39cc50513, /*  359 */
128'hd51783878713bfe99a8505130000d517, /*  360 */
128'hd51784078793fce608e39ba505130000, /*  361 */
128'h970505130000d517bf759ba505130000, /*  362 */
128'h84ae892af406e84aec26f02271798082, /*  363 */
128'h942a9041144201045513029044634401, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985ca808261459141694264e2, /*  366 */
128'h00f107a334f9090900c14783703050ef, /*  367 */
128'hbf55943e00e1578300f1072300d14783, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50563842e8067, /*  370 */
128'h082884b205e944079a638005079b0af5, /*  371 */
128'he517461985ca006409136b1050ef4611, /*  372 */
128'h07930174458369d050ef9d2505130000, /*  373 */
128'h1cf5826347b108b7e76332f5896302e0, /*  374 */
128'h478502b7e3631af58363479104b7e563, /*  375 */
128'h83638fa505130000d517478910f58463, /*  376 */
128'ha41d006040efa96505130000d51702f5, /*  377 */
128'h900505130000d51747a118f582634799, /*  378 */
128'h2cf5826347f5a4317ed030effef591e3, /*  379 */
128'h0000d51747d916f58a6347c500b7ed63, /*  380 */
128'h866302100793bf6dfef580e391c50513, /*  381 */
128'h05130000d517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5826306200793b7c99365, /*  383 */
128'h02f0079300b7ef632af5826303300793, /*  384 */
128'h938505130000d5170320079328f58763, /*  385 */
128'h079328f5846305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de394e505130000d51705e0, /*  387 */
128'h0670079300b7ef6328f5866308400793, /*  388 */
128'h960505130000d51706c0079326f58b63, /*  389 */
128'h079326f5886308900793b73df4f58ae3, /*  390 */
128'hd517f0f59ce30880079326f589630ff0, /*  391 */
128'h0000e79701e45703b73d96a505130000, /*  392 */
128'h12f714638dc989930000e9978e47d783, /*  393 */
128'h10f71c638ce7d7830000e79702045703, /*  394 */
128'h0000e597461953d050ef852285ca4619, /*  395 */
128'h012301a4578352d050ef854a89c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h0ea3db9ff0ef00f41e230029d78300f4, /*  399 */
128'h1223862601c1578300a10e23812100a1, /*  400 */
128'h0000c517a06ddcbfe0ef450185a202f4, /*  401 */
128'hb55977a505130000c517bd4176c50513, /*  402 */
128'h470302444783bdb5788505130000c517, /*  403 */
128'h178300f10e230254478300f10ea30264, /*  404 */
128'h00e10e2327810274470300e10ea301c1, /*  405 */
128'h0234470300e10ea301c1190302244703, /*  406 */
128'h04e79b6301c156830450071300e10e23, /*  407 */
128'h0000d597461947e27ad79e230000d797, /*  408 */
128'h0000d71779c505130000d51779458593, /*  409 */
128'hd79766a2476244d050efe43678f72e23, /*  410 */
128'h450102a40593ff89061b772787930000, /*  411 */
128'h616179a2794274e2640660a655e060ef, /*  412 */
128'h0000d71747e204e69463043007138082, /*  413 */
128'hc799439c760787930000d79774f72e23, /*  414 */
128'h0000d697f7e9439c750787930000d797, /*  415 */
128'h0000d597740606130000d61774468693, /*  416 */
128'h0713b765d6dfe0ef02a4051374458593, /*  417 */
128'h30ef6a2505130000c51702e798634d20, /*  418 */
128'h05130000c517cdcff0ef852285a65730, /*  419 */
128'hcc6ff0ef02a4051385ca55f030ef69e5, /*  420 */
128'h67c101e45703f6e787e35fe00713bf95, /*  421 */
128'h4611f4f70de302045703f6f701e317fd, /*  422 */
128'hb799379050ef0868700585930000d597, /*  423 */
128'h05130000c517b335678505130000c517, /*  424 */
128'hc517bb21694505130000c517b30d67e5, /*  425 */
128'h6b8505130000c517b3396a2505130000, /*  426 */
128'h0000c517b9ed6be505130000c517b311, /*  427 */
128'hb1dd6ea505130000c517b9c56dc50513, /*  428 */
128'h05130000c517b9f1700505130000c517, /*  429 */
128'hd703b1e1734505130000c517b9c97265, /*  430 */
128'h84930000d49767e7d7830000d7970265, /*  431 */
128'hd7830000d7970285d703ecf711e36764, /*  432 */
128'h89930205891320000793eaf719e36687, /*  433 */
128'h2c7050ef854a85ce461900f59a230165, /*  434 */
128'h2b7050ef854e626585930000d5974619, /*  435 */
128'h50ef00640513616585930000d5974619, /*  436 */
128'h01c4578329b050ef852285ca46192a50, /*  437 */
128'h02f4142301e4578302f4132302a00613, /*  438 */
128'h00f41f230024d78300f41e230004d783, /*  439 */
128'h0000c51785aab36900f4162360800793, /*  440 */
128'h430017b7bba5460140d030ef6bc50513, /*  441 */
128'h74132601608130239f0101138307b603, /*  442 */
128'h8406871b0387759366850034171b00f6, /*  443 */
128'h3c23630c8387b783972a430005379f2d, /*  444 */
128'h5f200813ffc5849b2581601134235e91, /*  445 */
128'h00c5963b101005938a1d08b8696335b9, /*  446 */
128'h87930000d797cfb527818ff1fff7c793, /*  447 */
128'h869b7007f7930084179bea25439054e7, /*  448 */
128'h00d100a3872646d496aa068e9ebd8006, /*  449 */
128'h00d100230086d69b0106d69b0106969b, /*  450 */
128'h806686936685c6918005069b00015503, /*  451 */
128'h67139fad377d8005859b658502d51a63, /*  452 */
128'h868a83f502d7473b1782270546a10077, /*  453 */
128'h862602e6446397c285b6430008378f95, /*  454 */
128'h30838287b823430017b70405aa1ff0ef, /*  455 */
128'h610101135f8134838526600134036081, /*  456 */
128'hbc2306a126050008380300d788338082, /*  457 */
128'he42643c0e8220c2007b71101b7e1ff06, /*  458 */
128'h16938304b703430014b747812401ec06, /*  459 */
128'h598505130000c517e7990206c1630337, /*  460 */
128'h64a2644260e2c3c00c2007b72d1030ef, /*  461 */
128'hf0227179bfc14785eb9ff0ef80826105, /*  462 */
128'h478585930000d597461184ae8432ec26, /*  463 */
128'h430787930000d7970ef050eff4060068, /*  464 */
128'h88930000d89785a6862247b20007a803, /*  465 */
128'hd5170450069341a757030000d7174168, /*  466 */
128'h740270a285228d4ff0ef422505130000, /*  467 */
128'h15428d5d05220085579b8082614564e2, /*  468 */
128'h8fd966c10185579b0185171b80829141, /*  469 */
128'h0085151b8fd98f750085571bf0068693, /*  470 */
128'h07b7715d808225018d5d8d7900ff0737, /*  471 */
128'h4581467d0390069300780207879b4b00, /*  472 */
128'hf052f44efc26e0a2f84ae486c63e4505, /*  473 */
128'h4d0505130000c517892a6ad070efec56, /*  474 */
128'h1d63c31901079713fff947931f1030ef, /*  475 */
128'hd717578538f706230000d71757b90a09, /*  476 */
128'h36f70d230000d717578938f701a30000, /*  477 */
128'h0000d717579136f708a30000d717578d, /*  478 */
128'hd797fe056513893d639070ef36f70423, /*  479 */
128'h34a585930000d597461134a78ba30000, /*  480 */
128'h338585930000d59746097e0050ef0048, /*  481 */
128'h06374722f2dff0ef45127d0050ef0028, /*  482 */
128'h77138ff183210087179bf00606130100, /*  483 */
128'hb02317c29101430016b78fd915020ff7, /*  484 */
128'h8086b7838006b78380f6b42393c180a6, /*  485 */
128'h79a2794274e282f6b42347a1640660a6, /*  486 */
128'h2d8484930000d497808261616ae27a02, /*  487 */
128'h863b4999404a0a130000ca175ae14401, /*  488 */
128'h56330286061b04852405855285a2028a, /*  489 */
128'h10e30f7030effec48fa30ff6761300c9, /*  490 */
128'h8087b5838007b603430017b7bf91ff34, /*  491 */
128'hf822fc068f4d91c115c2008007377139, /*  492 */
128'h80e7b423e05ae456e852ec4ef04af426, /*  493 */
128'h0000d7170b9030ef3c0505130000c517, /*  494 */
128'h0000d8172607c7830000d79726774703, /*  495 */
128'h0000d61724e6c6830000d69725984803, /*  496 */
128'h0000c51723c5c5830000d59724564603, /*  497 */
128'h228404130000d41707d030ef39450513, /*  498 */
128'hd717202989930000d997448100044783, /*  499 */
128'h0a130000da170014478320f70d230000, /*  500 */
128'h0024478320f702a30000d7176a891f6a, /*  501 */
128'h1ef709230000d7174300193700262b37, /*  502 */
128'h004447831ef703a30000d71700344783, /*  503 */
128'h0000d717005447831cf70e230000d717, /*  504 */
128'h0000d7971a0794230000d7971cf708a3, /*  505 */
128'h0000d7971a07a2230000d7971807ae23, /*  506 */
128'ha783e4a91807a6230000d7971807ac23, /*  507 */
128'h37835a0b0493ed9fe0ef8522e78d0009, /*  508 */
128'h97138309378302074563033797138309, /*  509 */
128'h000a2783bfc5bb7ff0effc075de30337, /*  510 */
128'hbfc1710a849377d050ef4501dff154fd, /*  511 */
128'h470300154783b7d914fdb7e9b9dff0ef, /*  512 */
128'h07c200354503002547838f5d07a20005, /*  513 */
128'h1363367d57fd808225018d5d05628fd9, /*  514 */
128'hfee50fa3058505050005c703808200f6, /*  515 */
128'h00b50023808200f61363367d57fdb7f5, /*  516 */
128'he04ae426ec06e8221101495cbfcd0505, /*  517 */
128'h02000513478101853903cfa500958413, /*  518 */
128'h0006c703462d02e0031348a5481586ca, /*  519 */
128'h95630e5007130107146300a70e632785, /*  520 */
128'h0685040500e400230405006400230117, /*  521 */
128'h842384ae01c9051300b94783fcc79ee3, /*  522 */
128'h0189470301994783c088f59ff0ef00f5, /*  523 */
128'h47030179478300f492238fd90087979b, /*  524 */
128'h0004002300f493238fd90087979b0169, /*  525 */
128'h873e611c80826105690264a2644260e2, /*  526 */
128'hfc630007468303a0061302000593cf99, /*  527 */
128'h577d00d706630017869300c6986302d5, /*  528 */
128'h869b577d46050007c683b7dd0705a00d, /*  529 */
128'h0006871b078900b666630ff6f593fd06, /*  530 */
128'hbfd5052747030000d7178082853ae11c, /*  531 */
128'h0067d683c70d0007c703cb85611cc915, /*  532 */
128'h0017c503e406114102e6906300855703, /*  533 */
128'h60a24525c3914501001577933f4060ef, /*  534 */
128'h01a5c70301b5c7838082452580820141, /*  535 */
128'h00d51d630007079b8f5d0087979b468d, /*  536 */
128'h979b8fd50087979b0145c6830155c783, /*  537 */
128'hec26f02271798082853e27818fd90107, /*  538 */
128'h842a03450993e052e84af4065904e44e, /*  539 */
128'h2501382060ef85ce8626468500154503, /*  540 */
128'heb6340f487bb000402234c58505ce131, /*  541 */
128'h6a0269a2694264e2740270a2450100e7, /*  542 */
128'h4c5cff2a74e34a050034490380826145, /*  543 */
128'h340060ef85ce86269cbd468500144503, /*  544 */
128'hf06fc39900454783b7f94505b7e5397d, /*  545 */
128'he426ec06e8221101591c80824501f8df, /*  546 */
128'hfddff0ef892e84aa02b787634401e04a, /*  547 */
128'h8593864a46850014c503ec190005041b, /*  548 */
128'ha823597d4405c11925012c8060ef0344, /*  549 */
128'h80826105690264a2644260e285220324, /*  550 */
128'h0005022357fde04ae426ec06e8221101, /*  551 */
128'h23344783e52d2501fa3ff0ef842ad91c, /*  552 */
128'h0107979b8fd90087979b450923244703, /*  553 */
128'h051302f71f63a55707134107d79b776d, /*  554 */
128'h0913010005370005079bd59ff0ef06a4, /*  555 */
128'h45010127f7b31465049300544537fff5, /*  556 */
128'h75332501d33ff0ef0864051300978c63, /*  557 */
128'h690264a2644260e200a035338d050125, /*  558 */
128'he486f44ef84a715dbfcd450d80826105, /*  559 */
128'h89aa00053023e85aec56f052fc26e0a2, /*  560 */
128'h171302054e6347addd9ff0ef8932852e, /*  561 */
128'h84aa638097bae56787930000d7970035, /*  562 */
128'h4503cb85000447830089b023c01547b1, /*  563 */
128'h00090563e38d00157793212060ef0014, /*  564 */
128'h79a2794274e2640660a647a9c1118911, /*  565 */
128'h0ff4f51380826161853e6b426ae27a02, /*  566 */
128'h00157713124060ef00a400a300040023, /*  567 */
128'h85224581f569891100090463fb71478d, /*  568 */
128'h1fa40913848a04f51a634785ee1ff0ef, /*  569 */
128'h854ac7894501ffc9478389a623a40a13, /*  570 */
128'h14e30991094100a9a0232501c5bff0ef, /*  571 */
128'h000a876345090004aa8301048913ff2a, /*  572 */
128'hfe9915e30491c10de9dff0ef852285d6, /*  573 */
128'h04e34785470db7bd00e519634785470d, /*  574 */
128'h470304044783bfb947b5c1194a81f6e5, /*  575 */
128'h4107d79b0107979b8fd90087979b03f4, /*  576 */
128'h04a4478304b44983fef711e320000713, /*  577 */
128'h490329811a09866300f9e9b30089999b, /*  578 */
128'h012401a3fff9079b470501342e230444, /*  579 */
128'h0164012304144b03faf769e30ff7f793, /*  580 */
128'h4a03ffc900fb77b3fffb079bfa0b03e3, /*  581 */
128'h142300fa6a33008a1a1b045447830464, /*  582 */
128'h0474448304844503f3c100fa77930144, /*  583 */
128'h47030434478314050e638d450085151b, /*  584 */
128'h033906bbdfb18fd90087979b25010424, /*  585 */
128'h64e3873200d7063b9f3d004a571b2781, /*  586 */
128'h6905dd8d84ae0364d5bb40c504bbf4c5, /*  587 */
128'h00b673630905165500b9393366411955, /*  588 */
128'hcc04d458015787bb248900ea873b490d, /*  589 */
128'hf00a15e310e91263470dd05c03542023, /*  590 */
128'h849b0024949bd408b17ff0ef06040513, /*  591 */
128'hc81c57fdee99e7e324810094d49b1ff4, /*  592 */
128'h08f91963478d00f402a3f8000793c45c, /*  593 */
128'h979b8fd90087979b0644470306544783, /*  594 */
128'h001a859b06f71b6347054107d79b0107, /*  595 */
128'h470323344783e13d2501ce5ff0ef8522, /*  596 */
128'h0107979b8fd90087979b000402a32324, /*  597 */
128'h051304f71263a55707134107d79b776d, /*  598 */
128'h252787932501416157b7a99ff0ef0344, /*  599 */
128'h614177b7a83ff0ef2184051302f51763, /*  600 */
128'hf0ef21c4051300f51c63272787932501, /*  601 */
128'hd797c448a63ff0ef22040513c808a6df, /*  602 */
128'h0000d71793c117c22785bdc7d7830000, /*  603 */
128'h00042a230124002300f41323bcf71723, /*  604 */
128'h0005099ba33ff0ef05840513b3514781, /*  605 */
128'he00a05e3b545a25ff0ef05440513b5b9, /*  606 */
128'hb7010014949b00f915634789d41c9fb5, /*  607 */
128'hbdc59cbd0017d79b8885029787bb478d, /*  608 */
128'h2501bffff0ef842ae426ec06e8221101, /*  609 */
128'h005447030cf71063478d00044703ed69, /*  610 */
128'h458120000613034404930af71b634785, /*  611 */
128'h079322f4092305500793a01ff0ef8526, /*  612 */
128'h0aa302f40a230520079322f409a3faa0, /*  613 */
128'h481c20f40da302f40b230610079302f4, /*  614 */
128'h0107971b20e40d2302e40ba304100713, /*  615 */
128'h20e40ea320f40e230087571b0107571b, /*  616 */
128'h0f23445c20f40fa30187d79b0107d71b, /*  617 */
128'h0087571b0107571b0107971b501020e4, /*  618 */
128'h22e400a322f400230720069300144503, /*  619 */
128'h0ca320d40c230187d79b0107d71b2605, /*  620 */
128'h85a64685d81022f401a322e4012320d4, /*  621 */
128'h4581460100144503000402a366d050ef, /*  622 */
128'h64a2644260e200a035332501661050ef, /*  623 */
128'h00f6f96337f9ffe5869b4d1c80826105, /*  624 */
128'h450180829d2d02d585bb554800254583, /*  625 */
128'hf406e84a71794d180eb7f76347858082, /*  626 */
128'h0005470302e5f963892ae44eec26f022, /*  627 */
128'h1e6308d70e63468d06d70c63842e4689, /*  628 */
128'h9dbd0094d59b9cad515c0015d49b00f7, /*  629 */
128'h64e2740270a257fdc9112501ac7ff0ef, /*  630 */
128'h899b0249278380826145853e69a26942, /*  631 */
128'h854a9dbd94ca1ff4f4930099d59b0014, /*  632 */
128'h1ff9f993f5792501a93ff0ef0344c483, /*  633 */
128'hc0198fc50087979b880503494783994e, /*  634 */
128'hd59b515cbf458fe9157d6505bf658391, /*  635 */
128'h0014141bfd592501a63ff0ef9dbd0085, /*  636 */
128'h979b034945030359478399221fe47413, /*  637 */
128'hf0ef9dbd0075d59b515cb7598fc90087, /*  638 */
128'h05131fc575130024151bf9352501a39f, /*  639 */
128'h17fd2501100007b7807ff0ef954a0345, /*  640 */
128'hf04a4540f82271398082853e4785b765, /*  641 */
128'h478500b51523e456e852ec4ef426fc06, /*  642 */
128'h790274a2744270e2450900f41c63892a, /*  643 */
128'h74e34f98611c808261216aa26a4269e2, /*  644 */
128'h00e69463470d0007c683e02184aefee4, /*  645 */
128'h28235788fce4f7e30087d703eb155798, /*  646 */
128'h88bd000937839d3d0044d79bd1710089, /*  647 */
128'h00993c2300a92a2394be034787930496, /*  648 */
128'h09925a7d843a0027c9838722b75d4501, /*  649 */
128'he59ff0ef0134f66385a2000935034a85, /*  650 */
128'h01440c630005041be6fff0efbf752501, /*  651 */
128'h84bbf6f476e34f9c00093783f68afbe3, /*  652 */
128'he822110100a55583b78d4505bfc14134, /*  653 */
128'he4950005049bf33ff0ef842aec06e426, /*  654 */
128'h6c08ec990005049b933ff0ef6008484c, /*  655 */
128'h802357156c1cf3cff0ef458102000613, /*  656 */
128'h8526644260e200e782234705601c00e7, /*  657 */
128'hf426f822fc06e85271398082610564a2, /*  658 */
128'h84aa4d1c16ba75634a05e456ec4ef04a, /*  659 */
128'h842e89324709000547830af5f0634989, /*  660 */
128'hda1b154794630ee78863470d0ae78f63, /*  661 */
128'hf0ef9dbd009a559b00ba0a3b515c0015, /*  662 */
128'h001a0a9b8805060996630005099b8b9f, /*  663 */
128'hc783014487b3cc191ffa7a130ff97793, /*  664 */
128'h8ff50049179b00f7f71316c166850347, /*  665 */
128'h8223478502fa0a239a260ff7f7938fd9, /*  666 */
128'h86bff0ef9dbd8526009ad59b50dc00f4, /*  667 */
128'h591bc40d1ffafa9300099f630005099b, /*  668 */
128'h82234785032a8a239aa60ff979130049, /*  669 */
128'h6a4269e2790274a2854e744270e200f4, /*  670 */
128'h591b0347c783015487b3808261216aa2, /*  671 */
128'h515cb7e90127e9339bc100f979130089, /*  672 */
128'h92e30005099b811ff0ef9dbd0085d59b, /*  673 */
128'h03240a2394261fe474130014141bfc09, /*  674 */
128'h03240aa30089591b0109591b0109191b, /*  675 */
128'hf0ef9dbd0075d59b515cbf7901448223, /*  676 */
128'h74130024141bf80996e30005099bfd8f, /*  677 */
128'h2501da0ff0ef85569aa603440a931fc4, /*  678 */
128'h94260109179b012569338d71f0000637, /*  679 */
128'h00fa80a30087d79b03240a230107d79b, /*  680 */
128'h012a81a300fa81230189591b0109579b, /*  681 */
128'hf822fc06ec4ef4267139bf3d4989b745, /*  682 */
128'h00c52903e19d89ae84aae456e852f04a, /*  683 */
128'h5afd4a05844a04f977634d1c04090a63, /*  684 */
128'ha8214401052a606304f4636324054c9c, /*  685 */
128'h57fd0887f86347850005041bc43ff0ef, /*  686 */
128'h790274a2744270e28522547d00f41d63, /*  687 */
128'h7ee3894e4c9c808261216aa26a4269e2, /*  688 */
128'hf0ef852685a24409bf554905b7d5faf4, /*  689 */
128'h11e305450863fd5507e3c9012501c05f, /*  690 */
128'hf0ef852685a2167d10000637b76dfb24, /*  691 */
128'h577dc4c0489c02099063e9052501de9f, /*  692 */
128'h0017e7930054c783c89c37fdfae783e3, /*  693 */
128'hdbbff0ef852685ce8622bf4900f482a3, /*  694 */
128'h7139bfad4405f6f50fe34785dd612501, /*  695 */
128'h030917932905f822fc0600a55903f04a, /*  696 */
128'h70e24511eb9993c1e456e852ec4ef426, /*  697 */
128'h808261216aa26a4269e2790274a27442, /*  698 */
128'h00099d63842a8a2e00f97993d7ed495c, /*  699 */
128'h071b00855783e18dc85c61082785480c, /*  700 */
128'h8793012415230996601cfcf775e30009, /*  701 */
128'h5a9b00254783bf5d4501ec1c97ce0347, /*  702 */
128'hb27ff0effc0a9fe30157fab337fd0049, /*  703 */
128'h57fdbf4945090097e46347850005049b, /*  704 */
128'h06f4e0634d1c6008b761450500f49463, /*  705 */
128'h451d0005049be81ff0ef480cf60a0ee3, /*  706 */
128'h6008fcf48de357fdfcf48be34785d4bd, /*  707 */
128'h4581200006136008f5792501dd8ff0ef, /*  708 */
128'h855285a600043a03beeff0ef03450513, /*  709 */
128'h0025478360084a0502aa2823aa5ff0ef, /*  710 */
128'hc8046008d91c415787bb591c00faed63, /*  711 */
128'hf0ef01450223b7b9c848a83ff0ef85a6, /*  712 */
128'hdb1c27855b1c2a856018f1412501d1cf, /*  713 */
128'he852ec4ef04afc06f426f8227139b7e9, /*  714 */
128'h842e84aa02f007130005c783e05ae456, /*  715 */
128'ha62304050ce7906305c0071300e78663, /*  716 */
128'h02f00a130ae7fc6347fd000447030004, /*  717 */
128'h8263000447834b2102e0099305c00a93, /*  718 */
128'h02000593462d0204b9030d5780630d47, /*  719 */
128'h00230d37926300044783b40ff0ef854a, /*  720 */
128'h00a302e007930b379063001447830139, /*  721 */
128'h09479763470d1b378e630024478300f9, /*  722 */
128'hf0ef8526458100f905a302000793943a, /*  723 */
128'hcdaff0ef608848cc100510632501adbf, /*  724 */
128'h00b74783c7e5000747836c98e96d2501, /*  725 */
128'h07050cb78d6300b78593709cef918ba1, /*  726 */
128'h4581fed608e3fff7c683fff746030785, /*  727 */
128'hb791c55c4bdc611cbf75dfdff0ef8526, /*  728 */
128'h70e20004bc232501a85ff0ef85264581, /*  729 */
128'h61216b026aa26a4269e2790274a27442, /*  730 */
128'h0693f7578be3bf954709bf1d04058082, /*  731 */
128'h4681b7ad02400793943a12f6e0630200, /*  732 */
128'h0505a0d1486502000313478145a14701, /*  733 */
128'h0023954a9101020695130027e793a8dd, /*  734 */
128'h069300094503c6ed4711a06d268500e5, /*  735 */
128'h0165966300d90023469500d515630e50, /*  736 */
128'h946345850037f6930ff7f7930027979b, /*  737 */
128'h671300d7946346918bb10107671300b6, /*  738 */
128'h4701bdfd00e905a39432920116020087, /*  739 */
128'h18e34711c50500b7c783709c4511bf65, /*  740 */
128'h0004a623cb890207f7930047f713f4e5, /*  741 */
128'h4515fb0dbf154501e80703e30004bc23, /*  742 */
128'hdbe58bc100b5c7836c8cfbf58b91b73d, /*  743 */
128'h9a63bdb9c4c8af2ff0ef0007c503609c, /*  744 */
128'h873245ad46a10ff7f7930027979b0565, /*  745 */
128'h74e3000747039722930117020017061b, /*  746 */
128'hf263fd370ae3f95704e3f94706e3f4e3, /*  747 */
128'hb51700054c634185551b0187151b02b6, /*  748 */
128'h10e30008866300054883412505130000, /*  749 */
128'h7ae30ff57513fbf7051bbd6d4519f117, /*  750 */
128'h3701eea866e30ff57513f9f7051beea8, /*  751 */
128'hec26f0227179bdf90ff777130017e793, /*  752 */
128'h0e500913451184aef406842ae44ee84a, /*  753 */
128'hafaff0ef6008a0b1c90de199484c49bd, /*  754 */
128'h00b7c783c3210007c7036c1ce1292501, /*  755 */
128'h17e18bfd033780630327026303f7f793, /*  756 */
128'h64e2740270a2450100979a630017b793, /*  757 */
128'hc13ff0ef852245818082614569a26942, /*  758 */
128'h1101bfe54511b7cd00042a23d9452501, /*  759 */
128'h250188fff0ef842ae426ec06e8224581, /*  760 */
128'h2501a8cff0ef6008484c0e500493e50d, /*  761 */
128'h4585cb9900978d630007c7836c1ced09, /*  762 */
128'h00f513634791dd792501bcdff0ef8522, /*  763 */
128'he82211018082610564a2644260e2451d, /*  764 */
128'he49d0005049bfa9ff0ef842aec06e426, /*  765 */
128'h6c08e0850005049ba42ff0ef6008484c, /*  766 */
128'h462d6c08700c84cff0ef458102000613, /*  767 */
128'h644260e200e782234705601c82aff0ef, /*  768 */
128'h450900b7ed6347858082610564a28526, /*  769 */
128'h6a0269a2694264e2740270a245098082, /*  770 */
128'he84af406ec26f02271794d1c80826145, /*  771 */
128'h59fd4a05fcf5fde384ae842ae052e44e, /*  772 */
128'h091bec8ff0ef852285a600f4fa634c1c, /*  773 */
128'h0763fb490ce3bf754501000914630005, /*  774 */
128'hf15d25018afff0ef852285a646010339, /*  775 */
128'he79300544783c81c278501378a63481c, /*  776 */
128'hb7594505bf5d0009049b00f402a30017, /*  777 */
128'hf0eff42ee432e82efc061028ec2a7139, /*  778 */
128'h050e0c2787930000c7970405426383ef, /*  779 */
128'h676200070023c3196622631800a78733, /*  780 */
128'h4785cb114501e39897aa00070023c319, /*  781 */
128'h2501a0eff0ef0828080c460100f61863, /*  782 */
128'he506f8ca7175bfe5452d8082612170e2, /*  783 */
128'h4925e42ee8daecd6f0d2f4cefca6e122, /*  784 */
128'h002c8a7984aa89b20005302314050d63, /*  785 */
128'h65a2140910630005091b9d6ff0ef1028, /*  786 */
128'he11964062501b6dff0efe4be1028083c, /*  787 */
128'hc54dc3e101f9fa1301c9f7934519e011, /*  788 */
128'h6a132501e75ff0ef102800f516634791, /*  789 */
128'h07937aa2cfcd008a77936406e949008a, /*  790 */
128'h072300f40ca300f408a3021007130460, /*  791 */
128'h0ba300040b2300e40823000407a30004, /*  792 */
128'h0ea300040e23000405a300e40c230004, /*  793 */
128'h85a2000ac50300040fa300040f230004, /*  794 */
128'h0a2300040da300040d234785fc9fe0ef, /*  795 */
128'h8b6300fa82230005099b00040aa30004, /*  796 */
128'h2501e3fff0ef030aab03855685ce0409, /*  797 */
128'h83aff0ef0135262385da39fd7522e911, /*  798 */
128'he3d98bc500b44783a895892ac90d2501, /*  799 */
128'h4783f565a0854921f60981e30049f993, /*  800 */
128'h000984630029f993e72d0107f71300b4, /*  801 */
128'h79a2020a6a13c399008a7793e3ad8b85, /*  802 */
128'h85a3d09c01448523f4800309a78385a2, /*  803 */
128'h01c40513c8c8f33fe0ef0009c5030004, /*  804 */
128'hae230004a623c8880069d783dbbfe0ef, /*  805 */
128'h854a640a60aa00f494230134b0230004, /*  806 */
128'h808261496b466ae67a0679a6794674e6, /*  807 */
128'he8d2eccef8a27119b7d5491db7e54911, /*  808 */
128'hf466f862fc5ee0daf0caf4a6fc86e4d6, /*  809 */
128'h8ab6e4328a2e842a0006a023ec6ef06a, /*  810 */
128'h00b44783000998630005099be91fe0ef, /*  811 */
128'h74a6854e744670e60007899bc39d6622, /*  812 */
128'h7ca27c427be26b066aa66a4669e67906, /*  813 */
128'h89638b8500a44783808261096de27d02, /*  814 */
128'h7463893e40f907bb445c010429031607, /*  815 */
128'h5c7d03040b1320000b930006091b00f6, /*  816 */
128'h6008120790631ff777934458fa090ce3, /*  817 */
128'hfc930197fcb337fd0025478300975c9b, /*  818 */
128'h00a7ec6347854848eb11020c99630ffc, /*  819 */
128'hbd6ff0ef4c0cb741498900f405a34789, /*  820 */
128'h498500f405a3478501851763b7e52501, /*  821 */
128'hb98ff0ef856e4c0c00043d83cc08b7a5, /*  822 */
128'h00a6073b0099579b000c861bd5792501, /*  823 */
128'hf4639fb1002dc683c4b58d3a0007849b, /*  824 */
128'h85d2863a86a6001dc503419684bb00f6, /*  825 */
128'h0407f79300a44783f94d250117a050ef, /*  826 */
128'h0097951b0097fc6341a507bb4c48c385, /*  827 */
128'hc5ffe0ef955285da2000061391011502, /*  828 */
128'h093b445c9a3e9381020497930094949b, /*  829 */
128'h00faa0239fa5000aa783c45c9fa54099, /*  830 */
128'h0407f79300a4478304e601634c50b705, /*  831 */
128'h140050efe43a85da4685001dc503c38d, /*  832 */
128'h0523fbf7f793672200a44783f1392501, /*  833 */
128'h50ef85da0017c503863a4685601c00f4, /*  834 */
128'h0009049b444c01a42e23f11525010ec0, /*  835 */
128'h0007849b0127f46340bb87bb1ff5f593, /*  836 */
128'hbf9dbd1fe0ef855295a2862603058593, /*  837 */
128'hfc56e0d2e4cee8caf0a27159b59d499d, /*  838 */
128'he46ee86aec66f062f45ef85aeca6f486, /*  839 */
128'hcb5fe0ef8ab689328a2e842a0006a023, /*  840 */
128'h899bc39d00b44783000997630005099b, /*  841 */
128'h6a0669a6694664e6854e740670a60007, /*  842 */
128'h61656da26d426ce27c027ba27b427ae2, /*  843 */
128'h873b445c18078f638b8900a447838082, /*  844 */
128'h5c7d03040b1320000b9304f76c630127, /*  845 */
128'h6008140793631ff77793040904634458, /*  846 */
128'hfc930197fcb337fd0025478300975c9b, /*  847 */
128'h4705cb914581485cef01040c9a630ffc, /*  848 */
128'h4c0cb759498900f405a3478902e79863, /*  849 */
128'h6a634818445cf3fd0005079bd86ff0ef, /*  850 */
128'hb79500f405230207e79300a4478312f7, /*  851 */
128'h4858bf99498500f405a3478501879763, /*  852 */
128'hc38d0407f79300a44783c85ce311cc1c, /*  853 */
128'h7e1040ef85da0017c50346854c50601c, /*  854 */
128'h00f40523fbf7f79300a44783f9692501, /*  855 */
128'hd159250197cff0ef856e4c0c00043d83, /*  856 */
128'h0007849b00a6863b0099579b000c869b, /*  857 */
128'h04bb00f774639fb5002dc703c4b58d32, /*  858 */
128'h2501793040ef85d286a6001dc5034197, /*  859 */
128'h0097959b0297f26341a587bb4c4cf151, /*  860 */
128'ha4ffe0ef855a95d22000061391811582, /*  861 */
128'h0094949b00f40523fbf7f79300a44783, /*  862 */
128'h9fa54099093b445c9a3e938102049793, /*  863 */
128'h4c5cbdd100faa0239fa5000aa783c45c, /*  864 */
128'h001dc50300e7fa63445c481800c78e63, /*  865 */
128'h01a42e23fd0925016f7040ef85da4685, /*  866 */
128'hf46340ab87bb1ff575130009049b4448, /*  867 */
128'h952285d28626030505130007849b0127, /*  868 */
128'h00f405230407e79300a447839dbfe0ef, /*  869 */
128'he406e0221141bd2d499db5f9c81cbf41, /*  870 */
128'hf71300a44783e1752501acffe0ef842a, /*  871 */
128'h46854c50601cc3950407f793cf690207, /*  872 */
128'hed5525016b5040ef030405930017c503, /*  873 */
128'h6008500c00f40523fbf7f79300a44783, /*  874 */
128'h671300b7c703741ce15d2501b77fe0ef, /*  875 */
128'h0106d69b0107169b481800e785a30207, /*  876 */
128'h0107569b00d78ea300e78e230086d69b, /*  877 */
128'h8b23485800e78fa300d78f230187571b, /*  878 */
128'h571b0107169b00e78d2300078ba30007, /*  879 */
128'h0107571b0107171b00e78a2327010107, /*  880 */
128'h021007130106d69b00e78aa30087571b, /*  881 */
128'h00d78da3046007130086d69b00e78c23, /*  882 */
128'h00a44783000789a30007892300e78ca3, /*  883 */
128'h00f50223478500f40523fdf7f7936008, /*  884 */
128'h640260a24505ebbfe06f014160a26402, /*  885 */
128'heffff0ef842ae406e022114180820141, /*  886 */
128'h3023e11925019cbfe0ef8522e9012501, /*  887 */
128'h0028e42a110180820141640260a20004, /*  888 */
128'h87230000c79700054a6395bfe0efec06, /*  889 */
128'h7159bfe5452d8082610560e245019ea7, /*  890 */
128'he0efeca6f486f0a21028002c4601e42a, /*  891 */
128'he4be1028083c65a2ec190005041bb3bf, /*  892 */
128'h77a2e9916586e41d0005041bcd2ff0ef, /*  893 */
128'h8082616564e6740670a68522cbd85752, /*  894 */
128'he0ef0004c50374a2cb998bc100b5c783, /*  895 */
128'hbfd94415fcf41ee34791b7c5c8c897bf, /*  896 */
128'hf0d2f4cef8cae122e506e42afca67175, /*  897 */
128'hacdfe0ef1828002c460184ae00050023, /*  898 */
128'h4bdc597d842677e2ecbe081ce5292501, /*  899 */
128'h67a24501040a12634a16c2be02f00993, /*  900 */
128'h80230307071b936747030000c717e505, /*  901 */
128'h07130e94186300e780a303a0071300e7, /*  902 */
128'h640a60aa00078023078d00e7812302f0, /*  903 */
128'h18284585808261497a0679a6794674e6, /*  904 */
128'he6eff0ef18284581fd452501f89fe0ef, /*  905 */
128'h8cdfe0ef0007c50365c677e2f5552501, /*  906 */
128'h4581f9492501f63fe0ef18284581c2aa, /*  907 */
128'hc50365c677e2e1052501e48ff0ef1828, /*  908 */
128'h1828458101450e6325018a7fe0ef0007, /*  909 */
128'hf8e516e367a24711dd612501a9eff0ef, /*  910 */
128'h97134781f5cfe0ef1828100cb7594509, /*  911 */
128'h871beb05fc9747039736109493010207, /*  912 */
128'h86bb40f405bbfff7871b04e462630037, /*  913 */
128'h01271a6396b2920166a20206961300e5, /*  914 */
128'hb7c12785b7319c3d01368023fff7c793, /*  915 */
128'h377dfc964603962a1088920102071613, /*  916 */
128'h169367220789bddd4545b7e900c68023, /*  917 */
128'h8fa32405078500074703973692810204, /*  918 */
128'hf04af426f8227139b709fe9465e3fee7, /*  919 */
128'hfb4fe0ef84ae842ae456e852ec4efc06, /*  920 */
128'h891bcf8900b44783000917630005091b, /*  921 */
128'h6a4269e2790274a2854a744270e20007, /*  922 */
128'h00a44783009777634818808261216aa2, /*  923 */
128'h445ce4bd00042623445884bae3918b89, /*  924 */
128'h0207e79300a44783c81cfcf778e34818, /*  925 */
128'hd3e51ff7f793445c4481bf7d00f40523, /*  926 */
128'hf7930304099300a44783fc960ee34c50, /*  927 */
128'h40ef0017c50385ce4685601cc3850407, /*  928 */
128'h0523fbf7f79300a44783ed51250133f0, /*  929 */
128'h40ef85ce0017c50386264685601c00f4, /*  930 */
128'h002547836008bf59cc44ed3525012ed0, /*  931 */
128'h0336d6bbfff4869b377dc7290097999b, /*  932 */
128'h4c0c8ff9413007bb02c6ed630337563b, /*  933 */
128'h0499ea634a855a7dd1c19c9dc45c2781, /*  934 */
128'he0ef6008d7b51ff4f793c45c9fa5445c, /*  935 */
128'h484cbfb19ca90094d49bcd112501c87f, /*  936 */
128'h00f5976347850005059b814ff0efe595, /*  937 */
128'h00f5976357fdbded490900f405a34789, /*  938 */
128'hb765cc0cc84cb5ed490500f405a34785, /*  939 */
128'h059bfddfe0efcb818b89600800a44783, /*  940 */
128'h0005059bc4bfe0efbf6984cee5990005, /*  941 */
128'hfaf5fae34f9c601cfabafee3fd4588e3, /*  942 */
128'hb7bdc45c013787bb413484bbcc0c445c, /*  943 */
128'h002c4601842ac52de42ef822fc067139, /*  944 */
128'h852265a267e2e1152501fe6fe0ef0828, /*  945 */
128'h6c0ce529250197cff0eff01c101ce01c, /*  946 */
128'h000430234515e7898bc100b5c783cd99, /*  947 */
128'h67e2c448e30fe0ef0007c50367e2a02d, /*  948 */
128'hcbdfe0ef00f414230067d78385224581, /*  949 */
128'h6121744270e2f971fcf50be347912501, /*  950 */
128'h1141b7c1fcf501e34791bfdd45258082, /*  951 */
128'h3023e1192501dbafe0ef842ae406e022, /*  952 */
128'hec26f022717980820141640260a20004, /*  953 */
128'h0005049bd98fe0ef892e842af406e84a, /*  954 */
128'h049bc5ffe0ef8522458100091f63e889, /*  955 */
128'h8082614564e269428526740270a20005, /*  956 */
128'h47912501b32ff0ef8522458102243023, /*  957 */
128'hc68fe0ef852285ca00042a2302f51363, /*  958 */
128'h00f5166347912501f8bfe0ef85224581, /*  959 */
128'heca67159bf6584aad16dbf7d00042a23, /*  960 */
128'he0eff486f0a21028002c460184aee42a, /*  961 */
128'he4be1028083c65a2e00d0005041bedaf, /*  962 */
128'hc489cf816786e8010005041b872ff0ef, /*  963 */
128'h64e6740670a68522c10fe0ef102885a6, /*  964 */
128'hf85a8432f0a27159bfcd441980826165, /*  965 */
128'heca6f486e0d28522002c46018b2ee42a, /*  966 */
128'he7cfe0efec66f062f45efc56e4cee8ca, /*  967 */
128'h481c01842c836000000a1c6300050a1b, /*  968 */
128'h740670a600fb202302f76263ffec871b, /*  969 */
128'h7ba27b427ae26a0669a6694664e68552, /*  970 */
128'h9f63478500044b83808261656ce27c02, /*  971 */
128'he0ef852285ca4a8559fd4481490902fb, /*  972 */
128'h2485e11109550863093508632501a55f, /*  973 */
128'he793c80400544783fef963e329054c1c, /*  974 */
128'h0ab7504cb74d009b202300f402a30017, /*  975 */
128'h00099e631afd4c094481498149011000, /*  976 */
128'h85cee9212501d10fe0ef0015899b8522, /*  977 */
128'h00194783038b91632000099303440913, /*  978 */
128'h09092485e3918fd90087979b00094703, /*  979 */
128'he0efe02e854ab745fc0c94e33cfd39f9, /*  980 */
128'h09112485e1116582015575332501abcf, /*  981 */
128'hbfad8a2abfbd4a09b7494a05b7c539f1, /*  982 */
128'hbc4fe0ef842ae04aec06e426e8221101, /*  983 */
128'h0007849bcb9100b44783e4910005049b, /*  984 */
128'h47838082610564a269028526644260e2, /*  985 */
128'hfed772e348144458cf390027f71300a4, /*  986 */
128'h484cef01600800f40523c8180207e793, /*  987 */
128'h00a405a3c53900042a232501a58ff0ef, /*  988 */
128'h57fd0005091b94dfe0ef4c0cbf7d84aa, /*  989 */
128'h167d100006374c0cb7dd450502f91463, /*  990 */
128'ha1cff0ef85ca6008f9792501b37fe0ef, /*  991 */
128'hfcf900e345094785b769449db7e12501, /*  992 */
128'h0407f79300a44783fcf96ae34d1c6008, /*  993 */
128'h030405930017c50346854c50601cdba5, /*  994 */
128'hfbf7f79300a44783f55d250171c040ef, /*  995 */
128'h1008002c4605e42a7175b7b100f40523, /*  996 */
128'he9052501ca0fe0eff8cafca6e122e506, /*  997 */
128'he1052501e3bfe0efe0be1008081c65a2, /*  998 */
128'h75e2eb890207f79300b7c78345196786, /*  999 */
128'h60aa451dcb810014f79300b5c483c599, /* 1000 */
128'h00094503790280826149794674e6640a, /* 1001 */
128'h2783c89d88c1cc0d0005041bad8fe0ef, /* 1002 */
128'he0ef00a8100c02800613fc878de30149, /* 1003 */
128'hf1612501951fe0efcaa200a8458996cf, /* 1004 */
128'h18e34791d94d2501836ff0ef00a84581, /* 1005 */
128'h7502e411f15525019f5fe0ef1008faf5, /* 1006 */
128'h91cff0ef85a27502bf612501f20fe0ef, /* 1007 */
128'h1028002c4605e42a7171b769d5752501, /* 1008 */
128'hf8dafcd6e152e54ee94aed26f506f122, /* 1009 */
128'h0005041bbd0fe0efe8eaece6f0e2f4de, /* 1010 */
128'hd67fe0efe4be1028083c65a21c041463, /* 1011 */
128'h67a61af4176347911c0409630005041b, /* 1012 */
128'h752218079f630207f79300b7c7834419, /* 1013 */
128'h4785180902630005091bb45fe0ef4581, /* 1014 */
128'h752216f90b63440557fd16f90f634409, /* 1015 */
128'h85ca7422160414630005041ba98fe0ef, /* 1016 */
128'h061303440a13f6efe0ef85220109549b, /* 1017 */
128'h462d898fe0ef855200050c1b45812000, /* 1018 */
128'hfb1347c1248188cfe0ef855202000593, /* 1019 */
128'hd99b02f40fa30104949b0109199b0ff4, /* 1020 */
128'h062302e00b930104d49b021007930109, /* 1021 */
128'hd49b0089d99b046007930ff97a9304f4, /* 1022 */
128'h052303740a230200061304f406a30084, /* 1023 */
128'h0423053407a305540723040405a30404, /* 1024 */
128'h80efe0ef0544051385d2049404a30564, /* 1025 */
128'h166357d200074603468d05740aa37722, /* 1026 */
128'h969b06f40723478100f69363571400d6, /* 1027 */
128'h0107979b06f4042327810107d79b0107, /* 1028 */
128'h0087d79b0086d69b0107d79b0106d69b, /* 1029 */
128'h99634c8500274b8306f404a306d407a3, /* 1030 */
128'h6786e8350005041bf59fe0ef1028040b, /* 1031 */
128'h00e78c230210071300e785a375224741, /* 1032 */
128'h00e78ca300078ba300078b2304600713, /* 1033 */
128'h00978aa301678a2301378da301578d23, /* 1034 */
128'ha82d0005041bd5afe0ef00f502234785, /* 1035 */
128'he0ef0195022303852823001c0d1b7522, /* 1036 */
128'h8552458120000613ec090005041b8dcf, /* 1037 */
128'h441db7498c6a0ffbfb93f61fd0ef3bfd, /* 1038 */
128'h64ea740a70aa8522f25fe0ef85ca7522, /* 1039 */
128'h6ce67c067ba67b467ae66a0a69aa694a, /* 1040 */
128'heca6f0a27159b7c544218082614d6d46, /* 1041 */
128'he0eff48610284605002c843284aee42a, /* 1042 */
128'he0efe4be1028083c65a2e13125019caf, /* 1043 */
128'hf79300b7c783451967a6e9152501b65f, /* 1044 */
128'h8cbd752200b74783c30d6706e39d0207, /* 1045 */
128'h02234785008705a38c3d027474138c65, /* 1046 */
128'h616564e6740670a62501c9efe0ef00f5, /* 1047 */
128'hf5060088002c4605e02ee42a71718082, /* 1048 */
128'h120796630005079b964fe0efed26f122, /* 1049 */
128'haf7fe0eff0be083cf4be008865a26786, /* 1050 */
128'h479900b7c703778610079a630005079b, /* 1051 */
128'h0e058e63479165e61007126302077713, /* 1052 */
128'h008c02800613e55fd0ef102805ad4655, /* 1053 */
128'h4d6347adf05fd0ef850ae49fd0ef10a8, /* 1054 */
128'hcbf90005079baadfe0ef10a865820c05, /* 1055 */
128'h0005079bdc5fe0ef10a80ce793634711, /* 1056 */
128'hd0ef00d4851302a10593464d648aefc5, /* 1057 */
128'h00f485a30207e793640602814783e0df, /* 1058 */
128'h4736cbbd8bc100b4c78300f402234785, /* 1059 */
128'hf2dfd0ef85a60004450306f7086357d6, /* 1060 */
128'h47890005059bcaefe0ef85220005059b, /* 1061 */
128'h6706efb10005079bfc3fd0ef8522c5a5, /* 1062 */
128'h969b57d602f69d630557468302e00793, /* 1063 */
128'h06f7042327810107d79b06f707230107, /* 1064 */
128'h0106d69b0087d79b0107d79b0107979b, /* 1065 */
128'h022306d707a3478506f704a30086d69b, /* 1066 */
128'h6506e7910005079be24fe0ef008800f7, /* 1067 */
128'h853e64ea740a70aa0005079bb50fe0ef, /* 1068 */
128'h842ee42ae8a2711dbfcd47a18082614d, /* 1069 */
128'he9292501810fe0efec861028002c4605, /* 1070 */
128'he12925019abfe0efe4be1028083c65a2, /* 1071 */
128'h6786eb950207f79300b7c783451967a6, /* 1072 */
128'h0087571b00e78b23752200645703cb85, /* 1073 */
128'h0087571b00e78c230044570300e78ba3, /* 1074 */
128'h2501ad6fe0ef00f50223478500e78ca3, /* 1075 */
128'he42ae0cae4a6711d80826125644660e6, /* 1076 */
128'hd0efec86e8a208284601002c893284ae, /* 1077 */
128'hd20208284581c4b9e0510005041bf9bf, /* 1078 */
128'hb8ffe0ef08284585e5592501ca8fe0ef, /* 1079 */
128'h8713ca1fd0ef8526462d75c2e93d2501, /* 1080 */
128'h879bce89000700230200061346ad00b4, /* 1081 */
128'h0007c78397a6938117820007869bfff6, /* 1082 */
128'hd0ef510c656202090a63fec783e3177d, /* 1083 */
128'h04300793470d6562e0150005041be69f, /* 1084 */
128'h034787930270079300e6846300054683, /* 1085 */
128'h644660e6852200a92023c29fd0ef953e, /* 1086 */
128'h802300f51563479180826125690664a6, /* 1087 */
128'h002c4605e42a711db7d5842abf550004, /* 1088 */
128'hec550005041bee3fd0efec86e8a21028, /* 1089 */
128'h97b6938102061793460100010c2366a2, /* 1090 */
128'h10284581ea2902000593eba10007c783, /* 1091 */
128'h10284585e8410005041bbd6fe0efda02, /* 1092 */
128'hc3dd650601814783e1792501abbfe0ef, /* 1093 */
128'h8c23021007136786bc7fd0ef082c462d, /* 1094 */
128'h8ca300078ba300078b230460071300e7, /* 1095 */
128'hfff6079bbf45863eb74d2605a06100e7, /* 1096 */
128'hfeb706e3000747039736930102079713, /* 1097 */
128'hc70348b107f00e9343658e2e4781082c, /* 1098 */
128'h00a36c6391411542f9f7051b27850006, /* 1099 */
128'h0f1be2a505130000a517934117423701, /* 1100 */
128'h644660e68522441900eef863a8210007, /* 1101 */
128'h0563000548030505bfcdf36d80826125, /* 1102 */
128'h00c6802300fe06b3b7cdffe81be30608, /* 1103 */
128'h02234785752200f500235795a8850785, /* 1104 */
128'h1b634791b7c10005041b8fefe0ef00f5, /* 1105 */
128'h041ba55fe0ef1028dbd50181478302f5, /* 1106 */
128'hb07fd0ef4581020006136506f4450005, /* 1107 */
128'h85a347216786ae5fd0ef082c462d6506, /* 1108 */
128'h00e58023f91780e3b751842abf1900e7, /* 1109 */
128'h0613472993811782f4c7e5e305850685, /* 1110 */
128'h079301814703f8d771e30007869b0200, /* 1111 */
128'h05452e0305052e83bf89eaf71de30e50, /* 1112 */
128'he44ae826ec22110105c5288305852303, /* 1113 */
128'h6f97887687f2869a8646040502938f2a, /* 1114 */
128'h00b647338dfd00c6c5b3a52f8f930000, /* 1115 */
128'h85bb0fc1008fa403000f2583000fa383, /* 1116 */
128'h0105883b004f2703ff4fa3839db90075, /* 1117 */
128'h0077073b0105e8330198581b0078159b, /* 1118 */
128'h23838e358e6d00f6c6339f3100f805bb, /* 1119 */
128'h83bb8e590146561b00c6171b9e39008f, /* 1120 */
128'h8ef900b7c6b300d383bb00c5873b0083, /* 1121 */
128'h969b00f6d39b007686bb8ebd00cf2403, /* 1122 */
128'h00d703bbffcfa4039fa100d3e6b30116, /* 1123 */
128'h9f3d8f2d9fa1007777338f2d0007061b, /* 1124 */
128'h0005881b0f418f5d0167171b00a7579b, /* 1125 */
128'h00006597f45f17e300e387bb0003869b, /* 1126 */
128'h000062979ccf8f9300006f97a9458593, /* 1127 */
128'h01e6c73300cf7f3300d7cf33a9428293, /* 1128 */
128'h00ef0f3b0025c4030015c383000faf03, /* 1129 */
128'h040a4318972a070a93aa038a0005c703, /* 1130 */
128'h1f1b010f083b004fa70300ef0f3b942a, /* 1131 */
128'h010f68330003a70301b8581b9e390058, /* 1132 */
128'h9e398e3d8e7501e7c6339f3100f80f3b, /* 1133 */
128'h40189eb90176561b0096139b008fa703, /* 1134 */
128'h007f46b305919f3500cf03bb00c3e633, /* 1135 */
128'ha7039eb90fc101e6c6b3fff5c4838efd, /* 1136 */
128'h0126d69b9fb900e6941b94aa048affcf, /* 1137 */
128'h77330083c7339fb900d3843b8ec14098, /* 1138 */
128'h0147171b00c7579b9f3d0077473301e7, /* 1139 */
128'h07bb0004069b0003861b000f081b8f5d, /* 1140 */
128'h8ffa9aaf0f1300006f17f25599e300e4, /* 1141 */
128'h0003a703010fc4039203839300006397, /* 1142 */
128'h9f25400000c2c4b3942a040a00d7c2b3, /* 1143 */
128'h9e2194aa048a0043a4039f21011fc483, /* 1144 */
128'h581b0048171b012fc4830107083b4080, /* 1145 */
128'h00f8073b0083a4039e210107683301c8, /* 1146 */
128'h408000c2863b9ea194aa00e2c2b3048a, /* 1147 */
128'h00c2e6330156561b013fc90300b6129b, /* 1148 */
128'h00e7c6b3ffc3a4839c3500c702bb03c1, /* 1149 */
128'h9fa50106941b992a9ea1090a0056c6b3, /* 1150 */
128'h081b00d2843b8ec1000924830106d69b, /* 1151 */
128'h0097579b9f3d8f219fa5005747330007, /* 1152 */
128'h0004069b0002861b0f918f5d0177171b, /* 1153 */
128'h8982829300006297f5f592e300e407bb, /* 1154 */
128'h43830002a70300d745b38f5dfff64713, /* 1155 */
128'h93aa038a020f45839f2d022f4403021f, /* 1156 */
128'h0042a5839f2d942a040a418c95aa058a, /* 1157 */
128'h581b0003a5839e2d0068171b0107083b, /* 1158 */
128'hfff6c6139db100f8073b0107683301a8, /* 1159 */
128'h561b00a6139b0082a5839e2d8e3d8e59, /* 1160 */
128'h9ead00c703bb00c3e633400c9ead0166, /* 1161 */
128'h8db902c10075e5b3fff7c593023f4483, /* 1162 */
128'hd59b94aa00f5969b048a9db5ffc2a403, /* 1163 */
128'h0007081b00b385bb40809fa18dd50115, /* 1164 */
128'h579b9f3d007747339fa18f4dfff74713, /* 1165 */
128'h869b0003861b0f118f5d0157171b00b7, /* 1166 */
128'h010e883b6462f3ef9de300e587bb0005, /* 1167 */
128'h0505282300c8863b00d306bb00fe07bb, /* 1168 */
128'h653c80826105692264c2cd70cd34c97c, /* 1169 */
128'he486e45ee85af44ef84afc26e0a2715d, /* 1170 */
128'h893289ae84aa97b203f7f413ec56f052, /* 1171 */
128'h8a1b408b07bb04000b9304000b13e53c, /* 1172 */
128'h1a9300090a1b00f97463938117820007, /* 1173 */
128'h043b86560084853385ce020ada93020a, /* 1174 */
128'h0174176399d641590933481020ef0144, /* 1175 */
128'h74e2640660a6b7c997824401852660bc, /* 1176 */
128'h808261616ba26b426ae27a0279a27942, /* 1177 */
128'he44eec26842a03f7f793f0227179653c, /* 1178 */
128'h802397a2f800071300178513e84af406, /* 1179 */
128'h0006091b40a9863b449d0400099300e7, /* 1180 */
128'h0124f5633c9020ef9522458192011602, /* 1181 */
128'hfde3450197828522603cfc1c078e643c, /* 1182 */
128'h8082614569a2694264e2740270a2fd24, /* 1183 */
128'he93c04053423639c4f0787930000a797, /* 1184 */
128'h00000797ed3c639c4e8787930000a797, /* 1185 */
128'h46410505059311018082e13cb6c78793, /* 1186 */
128'h86930000a69747013bf020efec06850a, /* 1187 */
128'h00e107b345418be585930000a5977566, /* 1188 */
128'h8bbd962e0047d613070506890007c783, /* 1189 */
128'h8fa3fec68f230007c78397ae00064603, /* 1190 */
128'h718505130000a51760e2fca71de3fef6, /* 1191 */
128'he42ee5060808842ae122717580826105, /* 1192 */
128'h0808e85ff0ef080885a26622f71ff0ef, /* 1193 */
128'h6149640a60aaf83ff0ef0808f01ff0ef, /* 1194 */
128'h1763469100d70d63711c46a159588082, /* 1195 */
128'h0007ac2380824501cf980200071300d7, /* 1196 */
128'h07b7ec06e426e82211018082556dbfe5, /* 1197 */
128'h86930000569702f5026384ae842a4200, /* 1198 */
128'ha517822585930000a597088006136466, /* 1199 */
128'h644260e2fc241cb030ef832505130000, /* 1200 */
128'hec06e4266100e82211018082610564a2, /* 1201 */
128'h86930000569702f4026384ae420007b7, /* 1202 */
128'h95177e2585930000959702f0061361e6, /* 1203 */
128'h644260e2e00418b030ef7f2505130000, /* 1204 */
128'hec06e4266100e82211018082610564a2, /* 1205 */
128'h86930000569702f4026384ae420007b7, /* 1206 */
128'h95177a25859300009597036006135ee6, /* 1207 */
128'h644260e2e40414b030ef7b2505130000, /* 1208 */
128'hec06e8226104e42611018082610564a2, /* 1209 */
128'h86930000a69702f48263842e420007b7, /* 1210 */
128'h9517762585930000959703e006134966, /* 1211 */
128'he8809001140210b030ef772505130000, /* 1212 */
128'h6104e42611018082610564a2644260e2, /* 1213 */
128'ha69702f48263842e420007b7ec06e822, /* 1214 */
128'h8593000095970450061344a686930000, /* 1215 */
128'h14020c7030ef72e505130000951771e5, /* 1216 */
128'h11018082610564a2644260e2ec809001, /* 1217 */
128'h026384ae420007b7ec06e4266100e822, /* 1218 */
128'h959704c00613536686930000569702f4, /* 1219 */
128'h30ef6ea50513000095176da585930000, /* 1220 */
128'h11018082610564a2644260e2f0040830, /* 1221 */
128'h026384ae420007b7ec06e4266100e822, /* 1222 */
128'h959705300613506686930000569702f4, /* 1223 */
128'h30ef6aa505130000951769a585930000, /* 1224 */
128'h71398082610564a2644260e2f4040430, /* 1225 */
128'h07b7fc06f04af426f82200053983ec4e, /* 1226 */
128'h0000569702f984638436893284ae4200, /* 1227 */
128'h650585930000959705a006134cc68693, /* 1228 */
128'h67227f6030efe43a6605051300009517, /* 1229 */
128'h004979130029191b8b0589890014159b, /* 1230 */
128'h744270e288a10125e5b30034949b8dd9, /* 1231 */
128'h8082612169e2790274a202b9b8238dc5, /* 1232 */
128'h458185224605468147057100e0221141, /* 1233 */
128'h8522f35ff0ef45818522f7dff0efe406, /* 1234 */
128'h45816008f67ff0ef4581460546854705, /* 1235 */
128'h1141808201414501640260a2d97ff0ef, /* 1236 */
128'h302302053c23460546814705e022e406, /* 1237 */
128'hf0ef45818522f39ff0ef842a45810405, /* 1238 */
128'hf23ff0ef46054685470545818522ef1f, /* 1239 */
128'h1101d4dff06f0141458160a264026008, /* 1240 */
128'h8263842e420007b7ec06e8226104e426, /* 1241 */
128'h9597061006133f6686930000569702f4, /* 1242 */
128'h30ef57a505130000951756a585930000, /* 1243 */
128'h610564a2644260e2fc80904114427120, /* 1244 */
128'h420007b7ec06e8226104e42611018082, /* 1245 */
128'h06133c2686930000569702f48263842e, /* 1246 */
128'h05130000951752658593000095970680, /* 1247 */
128'h60e2e0a08c7d17fd67856ce030ef5365, /* 1248 */
128'he4266100e82211018082610564a26442, /* 1249 */
128'h0000569702f4026384ae420007b7ec06, /* 1250 */
128'h4e0585930000959706f0061338c68693, /* 1251 */
128'h60e2e424688030ef4f05051300009517, /* 1252 */
128'h00053903e04a11018082610564a26442, /* 1253 */
128'h026384ae842a420007b7ec06e426e822, /* 1254 */
128'h959707600613356686930000569702f9, /* 1255 */
128'h30ef4aa505130000951749a585930000, /* 1256 */
128'h690264a2644260e2c84404993c236420, /* 1257 */
128'hf486e8caeca67100f0a2715980826105, /* 1258 */
128'h08a3ec66f062f45ef85afc56e0d2e4ce, /* 1259 */
128'h4611d01ce03084b2892e0005d7830204, /* 1260 */
128'h60080e049c636ca020ef00c905134581, /* 1261 */
128'h3a03420007b700043983bf5ff0ef4585, /* 1262 */
128'h0017f71344810049278316f99a630404, /* 1263 */
128'h03243c234c1c4485e391448d8b89c709, /* 1264 */
128'h160786638b85008a2783000a09638cdd, /* 1265 */
128'hf0ef852245814605468147050144e493, /* 1266 */
128'h852200892583be1ff0ef85224581d71f, /* 1267 */
128'h00095583c4fff0ef2d0c0c1300005c17, /* 1268 */
128'h85a6c81ff0ef3c6a0a1300009a178522, /* 1269 */
128'h4705cf5ff0ef85224581cbdff0ef8522, /* 1270 */
128'h000f45b7d27ff0ef8522458146054685, /* 1271 */
128'hf0ef85224585e93ff0ef852224058593, /* 1272 */
128'h0015e593009899b785220d89b583cd1f, /* 1273 */
128'h8a9300009a9768198993eb7ff0ef2581, /* 1274 */
128'h69a6694664e6740670a6efe9485c386a, /* 1275 */
128'h616545016ce27c027ba27b427ae26a06, /* 1276 */
128'h8522488cdb7ff0efe024852244cc8082, /* 1277 */
128'h3883603cee079be38b85449cdf3ff0ef, /* 1278 */
128'h47014781458163900107e68365410004, /* 1279 */
128'hec0689e36e89f005051300ff0e374311, /* 1280 */
128'he7b301e8183b070500371f1b00064803, /* 1281 */
128'hd81bf2e50067036316fd060527810107, /* 1282 */
128'h78330087981b010767330187971b0187, /* 1283 */
128'h873b8fd98fe9010767330087d79b01c8, /* 1284 */
128'h2585e31c9746938183751782170200be, /* 1285 */
128'h06131726869300005697b76547014781, /* 1286 */
128'h0513000095172a658593000095971490, /* 1287 */
128'h8b4ebd6100c4e493bd8544e030ef2b65, /* 1288 */
128'h859300005597000b1d633b7d42000bb7, /* 1289 */
128'hb7116f6000ef2a650513000095171565, /* 1290 */
128'h85d20f20061386e20179096300043903, /* 1291 */
128'h8cfd4c81485c0709348340e030ef8556, /* 1292 */
128'h6f630c8937830209370312048e632481, /* 1293 */
128'h85224581cc5cf9200793c7817c1c00f7, /* 1294 */
128'h0044f793b27ff0ef85224581b6fff0ef, /* 1295 */
128'h00896913ff397913852201442903c395, /* 1296 */
128'h248505130000951785cad47ff0ef85ca, /* 1297 */
128'h852201442903c3950084f793680000ef, /* 1298 */
128'h85cad1fff0ef85ca00496913ff397913, /* 1299 */
128'h0014f793658000ef2485051300009517, /* 1300 */
128'h5697017c8c630384390300043c83cfb5, /* 1301 */
128'h30ef855685d209c006130c2686930000, /* 1302 */
128'h470d02043c2300492783cba97c1c3620, /* 1303 */
128'h00c90793018c871308e69f630037f693, /* 1304 */
128'h0086161bff87051363104591480d4681, /* 1305 */
128'hc3988f518361ff87370301068763c390, /* 1306 */
128'h485ccbb5603cfeb690e30791872a2685, /* 1307 */
128'h4c858889c85c9bf9485cc85c0027e793, /* 1308 */
128'h0000569701748c63040439036004cc9d, /* 1309 */
128'h2e4030ef855685d20ca0061305c68693, /* 1310 */
128'hef8d8b85008927830009096304043023, /* 1311 */
128'h484cc85c9bf54c85485cb4dff0ef8522, /* 1312 */
128'h641020ef4505d80c8ee3c47ff0ef8522, /* 1313 */
128'hb77100f92623000cb783dbd98b85bd95, /* 1314 */
128'h0109648397a667a1bf41b1dff0ef8522, /* 1315 */
128'h639c00878913fa978de394be00093c83, /* 1316 */
128'h87ca0ca139a020efe43e002c46218566, /* 1317 */
128'hf02204800513717908b041635535b7dd, /* 1318 */
128'h1d4030ef892e84b2e44ef406e84aec26, /* 1319 */
128'hfc8505130000551785a2cc1d5551842a, /* 1320 */
128'h051300009517862285aa89aa785010ef, /* 1321 */
128'he01c420007b702098b634fe000ef1165, /* 1322 */
128'hc45c4789cb990024f793f40401242423, /* 1323 */
128'h8082614569a2694264e2740270a24501, /* 1324 */
128'h30ef8522b7e5c45c4785d4fd45018885, /* 1325 */
128'h42000537458146098082bff9557d1bc0, /* 1326 */
128'h25016108953e050e420007b7f73ff06f, /* 1327 */
128'h420007b7e4066380e0221141711c8082, /* 1328 */
128'h34c00613f64686930000569702f40263, /* 1329 */
128'h0085051300009517ff85859300009597, /* 1330 */
128'h640260a2557de3914505703c1a0030ef, /* 1331 */
128'he42eec064501842ae822110180820141, /* 1332 */
128'h6105468560e26622644285a24d3010ef, /* 1333 */
128'hec26f022f4062000051371797940006f, /* 1334 */
128'h0000951784aa0da030efe052e44ee84a, /* 1335 */
128'h44b010ef0001b5031e2030ef06c50513, /* 1336 */
128'h9517681c206010ef842a491010ef4501, /* 1337 */
128'h06f445833f8000ef638c052505130000, /* 1338 */
128'h9517546c3e8000ef0505051300009517, /* 1339 */
128'h00ef91c115c20085d59b05a505130000, /* 1340 */
128'h050505130000951706c44583583c3d20, /* 1341 */
128'h0ff777130187d61b0107d69b0087d71b, /* 1342 */
128'h5c0c3a6000ef26010ff6f6930ff7f793, /* 1343 */
128'h9597545c398000ef0405051300009517, /* 1344 */
128'hfb85859300009597c789fca585930000, /* 1345 */
128'h00009517378000ef0305051300009517, /* 1346 */
128'h8593000095977448132030ef03c50513, /* 1347 */
128'h00009617584c19c42783db7fb0ef6565, /* 1348 */
128'h95172f26061300009617e789f9460613, /* 1349 */
128'h84264581852633a000ef01a505130000, /* 1350 */
128'h999701aa0a1300009a174481ed5ff0ef, /* 1351 */
128'he78901f4f7932000091301a989930000, /* 1352 */
128'h2485854e0004458330c000ef855285a6, /* 1353 */
128'hfd249fe304052fa000ef819100f5f613, /* 1354 */
128'h740270a22e8000ef5e05051300009517, /* 1355 */
128'hb7038082614545016a0269a2694264e2, /* 1356 */
128'h278540f707b30003b6830083b7830103, /* 1357 */
128'h00f3b8230017079300d7fe6393811782, /* 1358 */
128'h80820007802345050103b78300a70023, /* 1359 */
128'h020596130103b7830083b70380824501, /* 1360 */
128'hf5638e9dfff706930003b7038f999201, /* 1361 */
128'hb70340a786bb87aa9d9dfff7059b00c6, /* 1362 */
128'h06938082852e0007002300b6e6630103, /* 1363 */
128'h00d7002307850007c68300d3b8230017, /* 1364 */
128'h488540a0053be681000556634881bfe9, /* 1365 */
128'h4e250ff6f81304100693c21906100693, /* 1366 */
128'h0ff3751302b6733b0005061b385986ba, /* 1367 */
128'h0ff5751302b6563b0305051b046e6763, /* 1368 */
128'h051340e685bbfe718532fea68fa30685, /* 1369 */
128'h802302d007930008876302f5e9630300, /* 1370 */
128'h000680230015559b40e6853b068500f6, /* 1371 */
128'h053b808200b61b63fff5081b86ba2581, /* 1372 */
128'h07bbb7d92585fea68fa30685bf5d00a8, /* 1373 */
128'h0006c8830007c30397ba9381178240c8, /* 1374 */
128'h7119b7f1068501178023006680232605, /* 1375 */
128'he4d6e8d2eccef4a6f8a2597d011cf0ca, /* 1376 */
128'hf82af02ef42afc3e843684b2e0dafc86, /* 1377 */
128'h0209591303000a9306c00a1302500993, /* 1378 */
128'h0017079bc52d8f1d0004c50377a27742, /* 1379 */
128'h04850135086304d7ff63938117827682, /* 1380 */
128'h0f630014c503bfe1e7bff0ef02010393, /* 1381 */
128'hcb9d0004c78303551063478104890545, /* 1382 */
128'h478100f6f36346a50ff7f793fd07879b, /* 1383 */
128'heb6306d50f630640069304890014c503, /* 1384 */
128'h09630630079304d50f630580069302a6, /* 1385 */
128'h6a4669e6790674a6744670e6f55d08f5, /* 1386 */
128'h0024c503808261090007051b6b066aa6, /* 1387 */
128'h00a76c6306e50e6307300713b74d048d, /* 1388 */
128'h4685003800840b13f6e51ee307000713, /* 1389 */
128'h0780071302e5006307500713a00d4601, /* 1390 */
128'h4685003800840b13fa850613f6e510e3, /* 1391 */
128'h00840b13f8b50693a81145c100163613, /* 1392 */
128'he37ff0ef400845a946010016b6930038, /* 1393 */
128'ha809ddbff0ef0028020103930005059b, /* 1394 */
128'hd93ff0ef00840b130201039300044503, /* 1395 */
128'h852201247433600000840b13b5fd845a, /* 1396 */
128'hb7f18522020103930005059b4db010ef, /* 1397 */
128'he4c6e0c2fc3ef83aec061034f436715d, /* 1398 */
128'hf032715d8082616160e2e8dff0efe436, /* 1399 */
128'hfc3ef83aec06100005931014862ef436, /* 1400 */
128'h8082616160e2e69ff0efe436e4c6e0c2, /* 1401 */
128'h100005931234862afe36fa32f62e710d, /* 1402 */
128'he436eec6eac2e6bee2baea22ee060808, /* 1403 */
128'h60f28522129020ef0808842ae3fff0ef, /* 1404 */
128'h03630087b303679c691c808261356452, /* 1405 */
128'h979304b7ee63479d8082450183020003, /* 1406 */
128'h439c97ba83f9abe70713000057170205, /* 1407 */
128'h2483795c878297bae426e822ec061101, /* 1408 */
128'h9381020497930c5010ef7540f55c08c5, /* 1409 */
128'h61054501e91c64a2644260e202f457b3, /* 1410 */
128'h058e05e135f1bfd9617cbfe97d5c8082, /* 1411 */
128'h11418082557d8082557db7e9659c95aa, /* 1412 */
128'h681c00055e63ff5ff0ef842ae406e022, /* 1413 */
128'h60a264028522000307630207b303679c, /* 1414 */
128'h557d80820141640260a2450183020141, /* 1415 */
128'h879300005797150200a7eb6347ad8082, /* 1416 */
128'h05130000951780826108953e8175a467, /* 1417 */
128'h715d83020007b303679c691c8082c165, /* 1418 */
128'h078517824785d23e47d502f1102347a1, /* 1419 */
128'hd402e486100c200007930030e83ee42e, /* 1420 */
128'h07374d148082616160a6fd3ff0efcc3e, /* 1421 */
128'h2381308345018082450100e6fe634004, /* 1422 */
128'h01138082240101132281348323013403, /* 1423 */
128'h342385a2980101f1041322813823dc01, /* 1424 */
128'hf579f95ff0ef1a05348322113c232291, /* 1425 */
128'h0dd4c70302f71c630a0447830a04c703, /* 1426 */
128'h0c0447830c04c70302f716630dd44783, /* 1427 */
128'h00f71a630e0447830e04c70302f71063, /* 1428 */
128'hd55156f010ef0d4485130d4405934611, /* 1429 */
128'h3e800513842af0227179b761fb600513, /* 1430 */
128'h00011023858a460185226ea020eff406, /* 1431 */
128'h7d000513e509842af21ff0efc202c402, /* 1432 */
128'h717980826145740270a285226cc020ef, /* 1433 */
128'hc402c23ef406f022478500f110234785, /* 1434 */
128'h87934ad4008007b745386914c195842a, /* 1435 */
128'h400006b78f75600006b78ff58ff9f807, /* 1436 */
128'hec9ff0ef8522858a4601c43e8fd98f55, /* 1437 */
128'h711d80826145740270a2c43c47b2e119, /* 1438 */
128'he0ca07c55783c23e47d500f1102347b5, /* 1439 */
128'h6a056989fdf949370107979bf852fc4e, /* 1440 */
128'h4495c43e842e8aaaec86f456e4a6e8a2, /* 1441 */
128'h858a4601e00a0a13e009899308090913, /* 1442 */
128'hc7891005f79345b2ed0de73ff0ef8556, /* 1443 */
128'h9517c78d0125f7b3054793630135f7b3, /* 1444 */
128'h60e6fba00513d4bff0efa72505130000, /* 1445 */
128'h808261257aa27a4279e2690664a66446, /* 1446 */
128'h00f057630014079b347dfe04c6e334fd, /* 1447 */
128'hfc8049e34501b7555d8020ef3e800513, /* 1448 */
128'hf9200513d09ff0efa485051300009517, /* 1449 */
128'h00f1102347c17139e7a919c52783bf7d, /* 1450 */
128'h842af426fc06f822858a460147d5c42e, /* 1451 */
128'hcb918b891b842783c11dde3ff0efc23e, /* 1452 */
128'h34fdc901dcdff0ef8522858a46014495, /* 1453 */
128'hbfd545018082612174a2744270e2f8ed, /* 1454 */
128'h4785e8a2ec86e0cae4a6711d80824501, /* 1455 */
128'h102302c9270347c906d7f66384b6892a, /* 1456 */
128'he42e4755d432cf3108c92783260102f1, /* 1457 */
128'hc83eca26d23a854a100c47850030cc3e, /* 1458 */
128'h47b10497f0634785e529842ad75ff0ef, /* 1459 */
128'hd23ed402854a100c47f5460102f11023, /* 1460 */
128'hf0ef9a25051300009517c11dd55ff0ef, /* 1461 */
128'h80826125690664a6644660e68522c43f, /* 1462 */
128'hb7d50004841bb74d02f6063bbf6147c5, /* 1463 */
128'hec4ef04af426f822fc067139b7c54401, /* 1464 */
128'h8ab684b28a2e4148842ace05e456e852, /* 1465 */
128'ha0ef852200b44583c11d892a482010ef, /* 1466 */
128'h00b67a63014485b3681000054d638c7f, /* 1467 */
128'ha0894481bd9ff0ef9585051300009517, /* 1468 */
128'h378389a6f96decdff0ef854a08c92583, /* 1469 */
128'h865286a2844e0089f3630207e4030109, /* 1470 */
128'h08c96783fc851ae3f01ff0ef854a85d6, /* 1471 */
128'hfc0999e39aa2028784339a22408989b3, /* 1472 */
128'h6aa26a4269e274a279028526744270e2, /* 1473 */
128'hc23e47f500f110234799713980826121, /* 1474 */
128'h8ed10106161b8edd030007b70086969b, /* 1475 */
128'h858a4601440dc43684aafc06f426f822, /* 1476 */
128'hf0ef85263e800593e919c53ff0ef8526, /* 1477 */
128'hfc79347d8082612174a2744270e2d91f, /* 1478 */
128'h23213823bffc07b7db0101134d18bfcd, /* 1479 */
128'h342322913c2324813023241134239fb9, /* 1480 */
128'h01f104131ce7f56349013ffc07372331, /* 1481 */
128'h1e051863892ac09ff0ef84aa85a29801, /* 1482 */
128'hb023796020ef20000513e7991a04b783, /* 1483 */
128'h85a2200006131e0503631a04b5031aa4, /* 1484 */
128'h47171cf76b6347210c044783123010ef, /* 1485 */
128'h400407b753b897ba078a5f2707130000, /* 1486 */
128'h67050d44278300e7fd63cc981ff78793, /* 1487 */
128'hf8dc00d773630147d69307a680070713, /* 1488 */
128'hf9938b8506f48f2309b449830a044783, /* 1489 */
128'h80a30b344783c7890e244783e7810019, /* 1490 */
128'h4783c7898b890a04478300098a6308f4, /* 1491 */
128'h8613091407130e24478306f48fa309c4, /* 1492 */
128'h468109d405130a844783fcdc07c60c84, /* 1493 */
128'h0087979b00074583fff74783e0fc07c6, /* 1494 */
128'h4685c39197aeffe745839fad0105959b, /* 1495 */
128'h0dd4478302f585b30e04458300098c63, /* 1496 */
128'hfca714e30621070de21c07ce02b787b3, /* 1497 */
128'h979b468508d4470308e4478304098f63, /* 1498 */
128'h470397ba08c447039fb90087171b0107, /* 1499 */
128'h07ce02e787b30dd4478302f707330e04, /* 1500 */
128'h171b0187979b08a4470308b44783f8fc, /* 1501 */
128'h47039fb90087171b089447039fb90107, /* 1502 */
128'h4783f4fc07a6c319f4fc54d89fb90884, /* 1503 */
128'hce81e3918bfd09c44783c7898b850a04, /* 1504 */
128'hed35e0bff0ef852645850af006134685, /* 1505 */
128'h8b850e0446830af447830af407a34785, /* 1506 */
128'h8663c79954dc08f4aa2300a6979bc7b9, /* 1507 */
128'h969b0dd44783f8dc07a60d4427830009, /* 1508 */
128'h80230a74478308d4ac2302f686bb00a6, /* 1509 */
128'h23813483854a240134032481308308f4, /* 1510 */
128'h50fc8082250101132281398323013903, /* 1511 */
128'h278527058bfd8b7d0057d79b00a7d71b, /* 1512 */
128'h1a04b503892abf4d08f4aa2302f707bb, /* 1513 */
128'hbf555951bf651a04b0235f8020efd169, /* 1514 */
128'h2281382322113c23dc010113bf455929, /* 1515 */
128'he16302f5886347892321302322913423, /* 1516 */
128'h230134032381308354a9c585468102b7, /* 1517 */
128'h80822401011322813483220139038526, /* 1518 */
128'h0613842e4685fef760e34705ffc5879b, /* 1519 */
128'h059bf57184aad1fff0ef892a45850b90, /* 1520 */
128'h85a2980101f10413f1e9258199f5ffe4, /* 1521 */
128'h0493f7d50b944783e51998dff0ef854a, /* 1522 */
128'he44ee84aec267179b74d84aab75ddf40, /* 1523 */
128'h0079f6930ff5f99308154783f022f406, /* 1524 */
128'hf0ef84aa45850b3006138edd892e9be1, /* 1525 */
128'h00091c6300f51e63842a57b5c519cc7f, /* 1526 */
128'h15e010ef8526842a875ff0ef852685ca, /* 1527 */
128'h69a2694264e2740270a28522013505a3, /* 1528 */
128'h2881382328113c23d601011380826145, /* 1529 */
128'h2741382327313c232921302328913423, /* 1530 */
128'h2581382325713c232761302327513423, /* 1531 */
128'he963478923b13c2325a1302325913423, /* 1532 */
128'h07b79f3dbff7879bbffc07b74d180ac7, /* 1533 */
128'h0000851784ae8b32892abfe787933ffc, /* 1534 */
128'h0016779307e9460300e7eb6355c50513, /* 1535 */
128'h0413f96ff0ef57e5051300008517e7b9, /* 1536 */
128'h2881348329013403298130838522f840, /* 1537 */
128'h26813a8327013a032781398328013903, /* 1538 */
128'h24813c8325013c0325813b8326013b03, /* 1539 */
128'h270380822a01011323813d8324013d03, /* 1540 */
128'h0045aa83db4555650513000085170989, /* 1541 */
128'hf7bb0005ac83e79102eaf7bb060a8163, /* 1542 */
128'hf24ff0ef55c5051300008517cb8902ec, /* 1543 */
128'he3994b8502eadabb02c92783bf415429, /* 1544 */
128'h478189d6856200c488138c0a009c9c9b, /* 1545 */
128'h02e8f33b0017859b000828834e114e85, /* 1546 */
128'hee4ff0ef554505130000851700030d63, /* 1547 */
128'h202302e8d33bb7f14b814a814c81b7c1, /* 1548 */
128'h8b850107c78397a6078e020880630065, /* 1549 */
128'h09bb0ffbfb9300dbebb300be96bbcb89, /* 1550 */
128'h000b8963fbc596e387ae051108210133, /* 1551 */
128'h0a13f00600e353650513000085178a09, /* 1552 */
128'h842af94ff0ef854a85d2fe0a7a1302f1, /* 1553 */
128'h0106161b09ea478309fa4603ee0519e3, /* 1554 */
128'h01367a63963e09da47839e3d0087979b, /* 1555 */
128'hb5c1e56ff0ef526505130000851785ce, /* 1556 */
128'hc71989b60017f7130a7a46830084c783, /* 1557 */
128'h450547010016e993c3990fe6f9938b89, /* 1558 */
128'h0017581b4b189726070e0017059b4611, /* 1559 */
128'h0027571b00b517bb0208046300187813, /* 1560 */
128'hd99b4187d79b8b050189999b0187979b, /* 1561 */
128'h92e3872e0ff9f99300f9e9b3c70d4189, /* 1562 */
128'h8517ef898b850a6a478302d98263fcc5, /* 1563 */
128'hfff7c793b5913a0020ef4da505130000, /* 1564 */
128'h8517cb898b8509ba4783bfd100f9f9b3, /* 1565 */
128'h02e3b51d547ddbaff0ef50a505130000, /* 1566 */
128'h0af006134685e3958b850afa4783e20b, /* 1567 */
128'h0afa07a34785e569a21ff0ef854a4585, /* 1568 */
128'h0880049308f92a2300a7979b0e0a4783, /* 1569 */
128'h86260ff6f69301acd6bb08c00d934d01, /* 1570 */
128'h0ff4f4932485ed499f1ff0ef854a4585, /* 1571 */
128'h019ad6bb08f00d134c81ffb492e32d21, /* 1572 */
128'he9359cbff0ef854a458586260ff6f693, /* 1573 */
128'h0d934d61ffa492e32ca10ff4f4932485, /* 1574 */
128'hd6bb45858656000c26834c818aa609b0, /* 1575 */
128'h2a85e13999dff0ef854a0ff6f6930196, /* 1576 */
128'h0ff4f493248dffac90e30ffafa932ca1, /* 1577 */
128'h854a458509c0061386defdb498e30c11, /* 1578 */
128'h0a7a4783d4fb0de34785ed19975ff0ef, /* 1579 */
128'hf0ef854a458509b00613468501379b63, /* 1580 */
128'h854a45850a70061386cebb3d842a957f, /* 1581 */
128'he406e0221141b32ddd79842a945ff0ef, /* 1582 */
128'hb303679c681c00055e63810ff0ef842a, /* 1583 */
128'h8302014160a264028522000307630187, /* 1584 */
128'hfc06f426713980820141640260a24505, /* 1585 */
128'h5529478500f5866384aa4791f04af822, /* 1586 */
128'h07c4d78300f110230370079304f59263, /* 1587 */
128'hc24a8526858a46010107979b4955842e, /* 1588 */
128'hc24a00f110234799ed19d52ff0efc43e, /* 1589 */
128'h8526858a4601c43e478900f41f634791, /* 1590 */
128'h80826121790274a2744270e2d34ff0ef, /* 1591 */
128'h4f5c6918ee09b7cdc402fef414e34785, /* 1592 */
128'h00e7f46385be27814f1887ae00f5f363, /* 1593 */
128'h8082c2cff06f02c50823dd0c0007059b, /* 1594 */
128'hf8a2070d4b9c711910000737691c8082, /* 1595 */
128'hfc5ee0dae4d6e8d2eccef0caf4a6fc86, /* 1596 */
128'hc509f11ff0ef842ac17c8fd9f466f862, /* 1597 */
128'h0000851702042423eb8d6b9c679c681c, /* 1598 */
128'h744670e6f8500493bacff0ef31c50513, /* 1599 */
128'h7be26b066aa66a4669e674a679068526, /* 1600 */
128'hf0eff3e54481541c808261097ca27c42, /* 1601 */
128'h2c2302f4082347851af42c23478df93f, /* 1602 */
128'h421010ef7d000513ba2ff0ef85220204, /* 1603 */
128'h2783f94584aa97826b9c679c8522681c, /* 1604 */
128'h478508f422231a04282318042e230884, /* 1605 */
128'hf0ef852245814601b72ff0ef8522d85c, /* 1606 */
128'h00ef8522f14984aacf2ff0ef8522f1df, /* 1607 */
128'h8737681c00f1102347a1000505a345d0, /* 1608 */
128'h0aa00713e3991aa007138ff94bdc00ff, /* 1609 */
128'hbf8ff0efc23ec43a8522858a460147d5, /* 1610 */
128'h07b700f715630aa0079300c14703e911, /* 1611 */
128'h0a934a55037009933e900913cc1c8002, /* 1612 */
128'h40000cb780020c3700ff8bb74b050290, /* 1613 */
128'hf0efc402c252013110238522858a4601, /* 1614 */
128'hc25a4bdc015110234c18681ce13dbb6f, /* 1615 */
128'hc43e0197e7b301871563c43e0177f7b3, /* 1616 */
128'hca6347b2ed1db8eff0ef8522858a4601, /* 1617 */
128'h331010ef3e80051306090863397d0007, /* 1618 */
128'h8001073700e68563800207374c14bf45, /* 1619 */
128'h06041e23d45c8b8541e7d79bc43ccc18, /* 1620 */
128'h02f51f63f9200793b55d18f40ca34785, /* 1621 */
128'hed09c34ff0ef85224581c04ff0ef8522, /* 1622 */
128'h4585bfd118f40c2347850007d663443c, /* 1623 */
128'h1985051300008517d965c1cff0ef8522, /* 1624 */
128'h551cb58584aab595fa100493a10ff0ef, /* 1625 */
128'hfed6e352e74eeb4aef26f706f3227161, /* 1626 */
128'he3b54401e6eeeaeaeee6f2e2f6defada, /* 1627 */
128'hc783c7b1199bc7831ff010ef45018baa, /* 1628 */
128'h460104f110234789e7b5180b8ca3198b, /* 1629 */
128'h842aabaff0efc482c2be855e008c479d, /* 1630 */
128'h46014495cf818b851b8ba783120500e3, /* 1631 */
128'h34fd100503e3842aaa0ff0ef855e008c, /* 1632 */
128'h842ad99ff0ef855ea031020ba423f4fd, /* 1633 */
128'h6a1a69ba695a64fa741a70ba8522d55d, /* 1634 */
128'h615d6db66d566cf67c167bb67b567af6, /* 1635 */
128'h855e0407c163180b8c23048ba7838082, /* 1636 */
128'h90810205149316d010ef4501b16ff0ef, /* 1637 */
128'hf155842ab36ff0ef855e45853e800913, /* 1638 */
128'h6ee3149010ef85260007cc63048ba783, /* 1639 */
128'h400007b7bfe91d7010ef0640051312a9, /* 1640 */
128'ha6238b8541e7d79b048ba78300fbac23, /* 1641 */
128'h1aa60f63450dbf0506fb9e23478502fb, /* 1642 */
128'h40010637a029400406370ea61ee34511, /* 1643 */
128'h49978a9d0036d61b00cbac234006061b, /* 1644 */
128'h460396ce964e068a8a3dc02989930000, /* 1645 */
128'h02d606bb018ba88345051086a6830f86, /* 1646 */
128'ha823180bae231a0ba8238a0500c7d61b, /* 1647 */
128'h8abd0107d69b08dba22308dba42304cb, /* 1648 */
128'h090ba8231408dc63090ba62300d5183b, /* 1649 */
128'h003f06b70107979b14068e6302cba683, /* 1650 */
128'h07854721938117828fd98ff50107571b, /* 1651 */
128'hb0230a0bbc23030787b300e797b30709, /* 1652 */
128'hb0230c0bbc230c0bb8230c0bb4230c0b, /* 1653 */
128'ha6230107d463200007930afbb8230e0b, /* 1654 */
128'ha82300e7f46320000793090ba70308fb, /* 1655 */
128'h471100e78e63577d04cba783c21508fb, /* 1656 */
128'hc4be04e11023855e008c46010107979b, /* 1657 */
128'h07cbd78304f11023479d902ff0efc282, /* 1658 */
128'hc4bec2ca855e008c0107979b46014955, /* 1659 */
128'h08fbaa234785e40516e3842a8e4ff0ef, /* 1660 */
128'h1ae3842ac9aff0ef855e08fb80a357fd, /* 1661 */
128'he0ef855e00b545830f7000ef855ee205, /* 1662 */
128'h54075a63018ba703e0051fe3842affbf, /* 1663 */
128'h10230370079304fba0232789100007b7, /* 1664 */
128'h855e0107979b108c460107cbd78306f1, /* 1665 */
128'h04934905d2caed05880ff0efd4bed2ca, /* 1666 */
128'h06f11023988102091a93033007930bf1, /* 1667 */
128'he826855e108c08104b210a854a11d482, /* 1668 */
128'hfe0a16e33a7dc131850ff0efd05aec56, /* 1669 */
128'hbd9940030637a7a940020637bb45842a, /* 1670 */
128'hb54d08bba82300b515bb89bd0165d59b, /* 1671 */
128'h8fd501e7569b8ff50027979b16f16685, /* 1672 */
128'h05374098b5558b1d938100f7571b1782, /* 1673 */
128'h8fd50087161b0187179b0187569b00ff, /* 1674 */
128'h8ef1f00706138fd167410087569b8e69, /* 1675 */
128'h169b0187559b40d804fbaa2327818fd5, /* 1676 */
128'h8ecd0087571b8de90087159b8ecd0187, /* 1677 */
128'h00638b3d0187d71b04ebac238f558f71, /* 1678 */
128'h00ebac238001073720d7026346892127, /* 1679 */
128'h20000737040ba7830007596302d79713, /* 1680 */
128'h1863800107b7018ba70304fba0238fd9, /* 1681 */
128'h040ba903639c5de78793000087971ef7, /* 1682 */
128'h00004497020d1a13044ba783f0be4d05, /* 1683 */
128'h83f979130ff1079300f97933a1c48493, /* 1684 */
128'h77b300e797bb478540980a05fe07fc13, /* 1685 */
128'h0b1b4a81017d8b3716078563278100f9, /* 1686 */
128'h00f977b340dc0007ac8397d6109c840b, /* 1687 */
128'h8d6345a1400007b7140781630197f7b3, /* 1688 */
128'h100005b700fc88634591200007b700fc, /* 1689 */
128'h8daa971ff0ef855e0015b59340bc85b3, /* 1690 */
128'h073700ec8d6347a1400007370e051c63, /* 1691 */
128'h40fc8cb3100007b700ec886347912000, /* 1692 */
128'h409cdfdfe0ef855e02fbaa23001cb793, /* 1693 */
128'h102347994d850ce79163470d01a78663, /* 1694 */
128'he7b317c12d81810007b7d33e47d50af1, /* 1695 */
128'he162855e110c040007930110d53e00fd, /* 1696 */
128'h8bbd010c4783e941e91fe0efc93ee552, /* 1697 */
128'ha58314079a631afba823409c09b79463, /* 1698 */
128'h18fbae2308bba2230017b79317ed088b, /* 1699 */
128'hfe07fd930ff10793947ff0ef855e4601, /* 1700 */
128'h4601475507cbd7830af1102303700793, /* 1701 */
128'hd53ee03ad33a8cee855e110c0107979b, /* 1702 */
128'hd33a0af1102347b56702e915e35fe0ef, /* 1703 */
128'he43e855e110c0110040007134791d502, /* 1704 */
128'h0e050c63e0dfe0efe03ac93ae552e16e, /* 1705 */
128'ha823017d85b74785f3ed37fd670267a2, /* 1706 */
128'h840585934601180bae23096ba2231afb, /* 1707 */
128'h04a1eafa94e347a10a918c9ff0ef855e, /* 1708 */
128'h00008517e6f49fe38987879300004797, /* 1709 */
128'h1737b61ddf400413cbdfe0efc7450513, /* 1710 */
128'h00ebac2380020737b519a007071b8001, /* 1711 */
128'h4905bbc580030737de075ee303079713, /* 1712 */
128'h3ac54a159881190201000ab70ff10493, /* 1713 */
128'h47d508f110234799020a08633a7d0905, /* 1714 */
128'hf426c556855e010c040007931030c33e, /* 1715 */
128'h83a54cdcd0051ce3d61fe0efdc3ef84a, /* 1716 */
128'h0087961bf006869366c144dcfbe18b85, /* 1717 */
128'h040ba70302e796938fd18ff50087d79b, /* 1718 */
128'h472db35d04fba02300876793da06d9e3, /* 1719 */
128'h2583974e837902079713eaf768e34581, /* 1720 */
128'h869300ff0537040d859366c1b5451187, /* 1721 */
128'h0187971b0187d61b0d91000da783f006, /* 1722 */
128'h8ff58f510087d79b8e690087961b8f51, /* 1723 */
128'h46a5008ca703fdb59ee3fefdae238fd9, /* 1724 */
128'h06b7018ba60300f6f8638bbd00c7579b, /* 1725 */
128'h078a6ea686930000369704d61c638003, /* 1726 */
128'ha68308fbae230087171b1487a78397b6, /* 1727 */
128'hd71b8fd10186d61b8ff917fd67c100cc, /* 1728 */
128'h3e800613c305c38d03f7771327810126, /* 1729 */
128'h06bb02f757bb8a8d0106d69b02e6073b, /* 1730 */
128'haa231b0ba7830adba2230afba02302d6, /* 1731 */
128'h08fba62320000793c79919cba7831afb, /* 1732 */
128'h062300051523484000ef855e08fba823, /* 1733 */
128'h8793ccccd6b7aaaab7b708cba7030005, /* 1734 */
128'h00d036b327818ef98ff9ccc68693aaa7, /* 1735 */
128'h0f068693f0f0f6b79fb500f037b30686, /* 1736 */
128'h8693ff0106b79fb5068a00d036b38ef9, /* 1737 */
128'h161376c19fb5068e00d036b38ef9f006, /* 1738 */
128'hb783d11c9fb9071200e037338f750207, /* 1739 */
128'hd68307abd70302c7d7b3ed1092010a8b, /* 1740 */
128'hab0585930000859784aa06fbc603074b, /* 1741 */
128'h070ba803a95fe0effef5362302450513, /* 1742 */
128'h0108571b0088579b06cbc603077bc883, /* 1743 */
128'h0ff777130ff878130ff7f7930188569b, /* 1744 */
128'he0ef04d48513a8e58593000085972681, /* 1745 */
128'h8513a8a5859300008597074ba603a5ff, /* 1746 */
128'he0ef8a3d8abd0146561b0106569b0624, /* 1747 */
128'hb8d102fba4234785015010ef8526a3ff, /* 1748 */
128'hb683400407b704fba0232785100007b7, /* 1749 */
128'ha085051300008517e691ecf76ce31a0b, /* 1750 */
128'hc78304fba0230017079b70000737bb95, /* 1751 */
128'hce910027f6931adba42303f7f6930c46, /* 1752 */
128'ha70304eba0230217071bc68900c7f693, /* 1753 */
128'ha783c7998b8504eba02301076713040b, /* 1754 */
128'ha783040baa0304fba02300c7e793040b, /* 1755 */
128'h349700fa7a33855e4601088ba583044b, /* 1756 */
128'h00003b174a85db4ff0ef59a484930000, /* 1757 */
128'h409c5dec8c9300003c974c2d5acb0b13, /* 1758 */
128'h00003917cbb5278100fa77b300fa97bb, /* 1759 */
128'h4703409c10000db720000d3758c90913, /* 1760 */
128'h270340dc04f718630017b79317ed0049, /* 1761 */
128'h061300894683c3a18ff900fa77b30009, /* 1762 */
128'hc131debfe0ef855e0fb6f69345850b70, /* 1763 */
128'ha783ddbfe0ef855e45850b7006134681, /* 1764 */
128'haa2308fba223180bae231a0ba823088b, /* 1765 */
128'h04a1fb9911e30931973fe0ef855e035b, /* 1766 */
128'h925fe0ef8dc5051300008517f7649fe3, /* 1767 */
128'h00d789634721400006b700092783bb6d, /* 1768 */
128'haa230017b71341b787b301a786634711, /* 1769 */
128'h808ff0ef855e408c933fe0ef855e02eb, /* 1770 */
128'ha823409ce79d0046f79300892683f941, /* 1771 */
128'ha2230017b79317ed088ba583ef8d1afb, /* 1772 */
128'h855ecb0ff0ef855e460118fbae2308bb, /* 1773 */
128'h0b7006130ff6f693bb91fd319fdfe0ef, /* 1774 */
128'h65e34581b7c9f521d31fe0ef855e4585, /* 1775 */
128'hbf6d11872583974e837902079713fcfc, /* 1776 */
128'h1023478d6da000ef06cb851300ec4641, /* 1777 */
128'hc4be0107979b008c460107cbd78304f1, /* 1778 */
128'hec051b63842a96ffe0efc2be47d5855e, /* 1779 */
128'h06fb9e2304e157830007d663018ba783, /* 1780 */
128'h460107cbd783c2be479d04f1102347a5, /* 1781 */
128'h842a93bfe0efc4be855e0107979b008c, /* 1782 */
128'h018ba50345e6475647c646b6ea051163, /* 1783 */
128'h06bba42306eba22306fba02304dbae23, /* 1784 */
128'h45098a3d01a6d61bf2c51a6340000637, /* 1785 */
128'h0637f0a609634505f0c543638ca602e3, /* 1786 */
128'hf06ffa100413f0eff06f2006061b4001, /* 1787 */
128'h8082557d8082557d80824501c56ce54f, /* 1788 */
128'h439c1de7879300008797808218b50d23, /* 1789 */
128'h00008717842ae406e02247851141ef9d, /* 1790 */
128'h5563aeefe0ef852212a000ef1cf72423, /* 1791 */
128'h13e000ef02c00513fc5ff0ef85220005, /* 1792 */
128'h4501808201414501640260a20dc000ef, /* 1793 */
128'h90636394631c19670713000087178082, /* 1794 */
128'he40688a505130000851785aa114102e7, /* 1795 */
128'ha60380820141853e478160a2f60fe0ef, /* 1796 */
128'h41488082853ebfd187b600a604630fc7, /* 1797 */
128'h10354703c105fbdff0efe42eec061101, /* 1798 */
128'h0c630ff007930815470302b7006365a2, /* 1799 */
128'h610560e25535eb3fe06f610560e200f7, /* 1800 */
128'he4261101bfcdf8400513bfe545018082, /* 1801 */
128'hf0ef842acd09f7dff0ef84aee822ec06, /* 1802 */
128'h64a2644260e2e0800f840413e501cf0f, /* 1803 */
128'hf807879300008797bfd5553580826105, /* 1804 */
128'h80820f8505138082c3980015071b4388, /* 1805 */
128'h8797110180824388f687879300008797, /* 1806 */
128'h84beec06e4266380e8220ca787930000, /* 1807 */
128'h47838082610564a2644260e200941763, /* 1808 */
128'h8797b7d56000a9cff0ef8522c78119a4, /* 1809 */
128'haf2300008797e79ce39c09a787930000, /* 1810 */
128'h67980827879300008797e5088082f007, /* 1811 */
128'h8497e4a6711d8082e308e518e11ce788, /* 1812 */
128'hf456f852fc4e6080e8a206a484930000, /* 1813 */
128'h89aae0caec86e06ae466e862ec5ef05a, /* 1814 */
128'h768a8a9300007a97778a0a1300007a17, /* 1815 */
128'h770b8b9300007b97770b0b1300007b17, /* 1816 */
128'h15634d29d54c8c9300007c9700050c1b, /* 1817 */
128'h7aa27a4279e2690664a660e664460294, /* 1818 */
128'h0513000085176d026ca26c426be27b02, /* 1819 */
128'h4c1cc7914901541cddcfe06f61258d65, /* 1820 */
128'h855a0fc42603681c89560007c3638952, /* 1821 */
128'he0ef855e85ca00090663dbefe0ef638c, /* 1822 */
128'hda4fe0ef856685e200978e63601cdb2f, /* 1823 */
128'h35a010efcdc505130000751701a98863, /* 1824 */
128'h4401e04ae426ec06e8221101b7716000, /* 1825 */
128'hcbad511ccbbd4d5ccfad44014d1cc141, /* 1826 */
128'h1c00059384aa892ec7ad639cc7bd651c, /* 1827 */
128'h4799c57c57fdcd21842a230010ef4505, /* 1828 */
128'h03253023e90410f502a347850ef52c23, /* 1829 */
128'h91c78793fffff797e65ff0ef04052823, /* 1830 */
128'h18f430232ee787930000179716f43c23, /* 1831 */
128'h2e23681c18f434232de7879300001797, /* 1832 */
128'he99ff0ef10f400230247c78385220ea4, /* 1833 */
128'h106f80826105690264a2644260e28522, /* 1834 */
128'h65186294611cc5668693000086971ec0, /* 1835 */
128'h0127d713e11897360017671302d786b3, /* 1836 */
128'h17bb40f007b300f7553b93ed836d8f3d, /* 1837 */
128'hee05051300008517808225018d5d00f7, /* 1838 */
128'h842afefff0efe022e4061141fc3ff06f, /* 1839 */
128'h2501640260a28d410105151bfe9ff0ef, /* 1840 */
128'h041bfdbff0efe022e406114180820141, /* 1841 */
128'h60a28d4115029001fd1ff0ef14020005, /* 1842 */
128'h0785fff5c703058587aa808201416402, /* 1843 */
128'h00c7896387aa962a8082fb75fee78fa3, /* 1844 */
128'h8082fb65fee78fa30785fff5c7030585, /* 1845 */
128'hc7030585eb09001786930007c70387aa, /* 1846 */
128'hb7d587b68082fb75fee78fa30785fff5, /* 1847 */
128'h001786930007c70387b68082e21987aa, /* 1848 */
128'h0fa300178713fff5c6830585963efb7d, /* 1849 */
128'h8082000780a300c715638082e291fed7, /* 1850 */
128'h07bbfff5c783000547030585b7cd87ba, /* 1851 */
128'hf37d0505e3994187d79b0187979b40f7, /* 1852 */
128'h0585a839478100c59463962e8082853e, /* 1853 */
128'h0187979b40f707bbfff5c78300054703, /* 1854 */
128'hf5938082853eff790505e3994187d79b, /* 1855 */
128'h0505c399808200b79363000547830ff5, /* 1856 */
128'h9363000547830ff5f59380824501bfcd, /* 1857 */
128'h0007c70387aabfcd0505dffd808200b7, /* 1858 */
128'he8221101bfcd0785808240a78533e701, /* 1859 */
128'hf593952265a2fe5ff0efec06842ae42e, /* 1860 */
128'hfe857be3157d00b78663000547830ff5, /* 1861 */
128'h856387aa95aa80826105644260e24501, /* 1862 */
128'h0785808240a78533e7010007c70300b7, /* 1863 */
128'hea9940c785330007c68387aa862ab7fd, /* 1864 */
128'hfe081be3000748030705fed80fe38082, /* 1865 */
128'h0007c60387aa86aabfcd872eb7d50785, /* 1866 */
128'h4803070500c80a638082ea1140d78533, /* 1867 */
128'hbff90785bfd5872e8082fe081be30007, /* 1868 */
128'h0785fee68fe380824501eb1900054703, /* 1869 */
128'h1101bfd587aeb7e50505fafd0007c683, /* 1870 */
128'h00008797e519842a84aeec06e426e822, /* 1871 */
128'hf9dff0ef85a68522cc116380cdc78793, /* 1872 */
128'hcc07b02300008797ef8100044783942a, /* 1873 */
128'h85a68082610564a2644260e285224401, /* 1874 */
128'h0023c78100054783c519f9fff0ef8522, /* 1875 */
128'h1101bfd9c8a7ba230000879705050005, /* 1876 */
128'hf0ef8526842ac891e822ec066104e426, /* 1877 */
128'h644260e2e008050500050023c501f73f, /* 1878 */
128'hcf9900054783c11d8082610564a28526, /* 1879 */
128'h8082e3110017c703ce810007c68387aa, /* 1880 */
128'h80824501b7e5078900d780a300e78023, /* 1881 */
128'h808204c79063963e87aacb9d00757793, /* 1882 */
128'h469d00c508b3872aff6d377d8fd507a2, /* 1883 */
128'h87335761003657930106ef6340e88833, /* 1884 */
128'h0ff5f6934725bfc1963a97aa078e02e7, /* 1885 */
128'hfeb78fa30785bfe1fef73c230721bfd1, /* 1886 */
128'h87aacb9d8b9d00a5e7b300b50a63bf6d, /* 1887 */
128'h07a1ff8738030721808202c79e63963e, /* 1888 */
128'h00365713ff06e8e340f88833ff07bc23, /* 1889 */
128'h00e507b3963e95ba070e02f707b357e1, /* 1890 */
128'h0585bfe1469d00c508b387aa872ebfc1, /* 1891 */
128'hf0227179bf65fee78fa30785fff5c703, /* 1892 */
128'hf0efe02ee84af406e432ec26852e842a, /* 1893 */
128'h00c564636582892ace1184aa6622dcdf, /* 1894 */
128'h0023f79ff0ef944a864a8522fff60913, /* 1895 */
128'h8082614564e269428526740270a20004, /* 1896 */
128'hf57ff0ef00a5e963842ae406e0221141, /* 1897 */
128'h00c506b395b280820141640260a28522, /* 1898 */
128'h0005c78315fdd7e500e587b340b60733, /* 1899 */
128'h478100c51563962ab7fd00f6802316fd, /* 1900 */
128'hfbed9f990005c703000547838082853e, /* 1901 */
128'h4783808200c51363962ab7dd05850505, /* 1902 */
128'h842af0227179bfc50505feb78de30005, /* 1903 */
128'hd1fff0ef89aee84af406e44eec26852e, /* 1904 */
128'h0005091bd13ff0ef8522c8890005049b, /* 1905 */
128'h694264e2740270a28522440100995b63, /* 1906 */
128'hf0ef397d852285ce86268082614569a2, /* 1907 */
128'h14630ff5f593962abfe90405d175f8bf, /* 1908 */
128'h0be300150793000547038082450100c5, /* 1909 */
128'h00c7ef630ff5f59347c1b7ed853efeb7, /* 1910 */
128'h0007c7038082853e4781e60187aa2601, /* 1911 */
128'hc31d00757713b7f5367d0785feb71ce3, /* 1912 */
128'h0007c80387aa0007069b40e7873b47a1, /* 1913 */
128'h938102071793faf5078536fdfcb81ce3, /* 1914 */
128'h0107179300b7e733008597938e1d953e, /* 1915 */
128'h87aa27018edd00365713020796938fd9, /* 1916 */
128'h0785f8b71fe30007c703d24d8a1deb11, /* 1917 */
128'h00d80a63008785130007b803bfcd367d, /* 1918 */
128'hbfa5fef51be30785f8b712e30007c703, /* 1919 */
128'h079300054703e7a9419cb7f1377d87aa, /* 1920 */
128'h8793000027970015470308f711630300, /* 1921 */
128'h071bc6898a850006c68300e786b36e67, /* 1922 */
128'h470304d71b63078006930ff777130207, /* 1923 */
128'h47c1c3b10447f7930007c78397ba0025, /* 1924 */
128'h07930005470302f71c6347c14198c19c, /* 1925 */
128'h0713000027170015478302f716630300, /* 1926 */
128'h0207879bc7098b0500074703973e6967, /* 1927 */
128'h8082050900e79363078007130ff7f793, /* 1928 */
128'h006c842ee8221101bf6d47a9bf7d47a1, /* 1929 */
128'h2817468100c16583f63ff0efc632ec06, /* 1930 */
128'h06330007079b00054703652808130000, /* 1931 */
128'hec0500089863044678930006460300f8, /* 1932 */
128'h8b6300467893808261058536644260e2, /* 1933 */
128'h050502d586b3feb7f4e3fd07879b0008, /* 1934 */
128'h0ff7f793fe07079bc6098a09b7d196be, /* 1935 */
128'hf426f8227139b7e1e008b7cdfc97879b, /* 1936 */
128'hf0ef84b2842ae42e00063023f04afc06, /* 1937 */
128'h790274a2744270e25529e90165a2b0df, /* 1938 */
128'hf5dff0ef8522082c892a862e80826121, /* 1939 */
128'h07858f81cb010007c703fe8782e367e2, /* 1940 */
128'hb7e94501e088fcf718e347a9fd279be3, /* 1941 */
128'hf2dff06f00e6846302d0071300054683, /* 1942 */
128'h40a0053360a2f23ff0efe40605051141, /* 1943 */
128'hf0dff0ef842ee406e022114180820141, /* 1944 */
128'hea6302d704630007c70304b00693601c, /* 1945 */
128'h0141640260a202d70e630470069300e6, /* 1946 */
128'h16e306b0069302d7076304d006938082, /* 1947 */
128'hfce69fe3052a069007130017c683fed7, /* 1948 */
128'he01c078d00e69863042007130027c683, /* 1949 */
128'he8221101bfd50789bff1052a052ab7e9, /* 1950 */
128'h00c16583e0fff0efc632ec06006c842e, /* 1951 */
128'h079b000547034fe80813000028174681, /* 1952 */
128'h9863044678930006460300f806330007, /* 1953 */
128'h7893808261058536644260e2ec050008, /* 1954 */
128'h86b3feb7f4e3fd07879b00088b630046, /* 1955 */
128'hfe07079bc6098a09b7d196be050502d5, /* 1956 */
128'h1141b7e1e008b7cdfc97879b0ff7f793, /* 1957 */
128'h04b00693601cf87ff0ef842ee406e022, /* 1958 */
128'h0470069300e6ea6302d704630007c703, /* 1959 */
128'h04d0069380820141640260a202d70e63, /* 1960 */
128'h0017c683fed716e306b0069302d70763, /* 1961 */
128'h07130027c683fce69fe3052a06900713, /* 1962 */
128'h052a052ab7e9e01c078d00e698630420, /* 1963 */
128'he589842ae406e0221141bfd50789bff1, /* 1964 */
128'h00002797fff5c70300a405b395bff0ef, /* 1965 */
128'h8b1100074703973efff5851342478793, /* 1966 */
128'h7ae3157d80820141557d640260a2e719, /* 1967 */
128'hf77d8b1100074703973e00054703fea4, /* 1968 */
128'hd7dff06f014105054581462960a26402, /* 1969 */
128'h0723812100a107a31141fa5ff06f4581, /* 1970 */
128'h8793000087978082014100e1550300a1, /* 1971 */
128'hf06f95be9201160291811582639c8b67, /* 1972 */
128'h853ee3190005470345a946254781aa5f, /* 1973 */
128'h87bb00d667630ff6f693fd07069b8082, /* 1974 */
128'he0221141bff90505fd07879b9fb902f5, /* 1975 */
128'h45a900b7f86347a500a04563842ee406, /* 1976 */
128'h02a4753b4529fe7ff0ef357d02b455bb, /* 1977 */
128'h07935000006f03050513014160a26402, /* 1978 */
128'h0000871782f73e230000871707e20810, /* 1979 */
128'h041300008417e8221101808282f73e23, /* 1980 */
128'hf0efec06600885aa84ae862ee42682e4, /* 1981 */
128'h610564a26442e00c95a660e2600ca15f, /* 1982 */
128'h7497e426804787930000879711018082, /* 1983 */
128'h000075176380e82260907f2484930000, /* 1984 */
128'h6088b87fd0ef85a29c11ec06cfc50513, /* 1985 */
128'h00007517862286aa608ce63fc0ef85a2, /* 1986 */
128'hd005051300007517b6dfd0efcf450513, /* 1987 */
128'h84bf90efef65051300000517b61fd0ef, /* 1988 */
128'h751740a005b364a260e2644200055e63, /* 1989 */
128'h60e26442b39fd06f6105cf2505130000, /* 1990 */
128'h8432e406e02211416980006f610564a2, /* 1991 */
128'h0141640260a2557d0085036386cfa0ef, /* 1992 */
128'he64e01258413f2227169808245018082, /* 1993 */
128'hf7eff0ef892eea4aee26f606852289aa, /* 1994 */
128'h95260505f72ff0ef852600a404b30505, /* 1995 */
128'h04e7ee631ff00793fff5071be93ff0ef, /* 1996 */
128'h84aaf50ff0ef852270a7ac2300007797, /* 1997 */
128'h07939526f42ff0efa685051300007517, /* 1998 */
128'h7517842af32ff0ef852204a7f2630ff0, /* 1999 */
128'h751700a405b3f24ff0efa4a505130000, /* 2000 */
128'h64f2741270b2a8bfd0efc62505130000, /* 2001 */
128'h00007717200007938082615569b26952, /* 2002 */
128'hf0ef850a458110000613b7556af72e23, /* 2003 */
128'hdeaff0ef850aa065859300007597863f, /* 2004 */
128'h0000759700f7096302f0079301294703, /* 2005 */
128'hf0ef850a85a2dfaff0ef850ac3458593, /* 2006 */
128'h7517858a43906767879300007797df2f, /* 2007 */
128'h07e208100793a1bfd0efc1a505130000, /* 2008 */
128'h3f230000771764f73f23000077174511, /* 2009 */
128'h450142a79d2300007797d85ff0ef64f7, /* 2010 */
128'h7597461142a7972300007797d77ff0ef, /* 2011 */
128'h77174785eb1ff0ef854e422585930000, /* 2012 */
128'he426ec06e8221101b79160f71f230000, /* 2013 */
128'h84ae450d892a08c7df638432478de04a, /* 2014 */
128'h751708a7956325010004d783d37ff0ef, /* 2015 */
128'h25010024d783d21ff0ef5ee555030000, /* 2016 */
128'hdabff0ef00448513ffc4059b06a79a63, /* 2017 */
128'h75173aa79d2300007797d05ff0ef4511, /* 2018 */
128'h000077974611cf1ff0ef5be555030000, /* 2019 */
128'hf0ef854a39c58593000075973aa79323, /* 2020 */
128'h5945d58300007597256000ef4535e2bf, /* 2021 */
128'h7797240000ef02000513d1bff0ef4515, /* 2022 */
128'h0000771727850007d78357e787930000, /* 2023 */
128'h278d439c564787930000779756f71823, /* 2024 */
128'h905fd0efb2450513000075170087cf63, /* 2025 */
128'h60e2d49ff06f6105690264a260e26442, /* 2026 */
128'hf022f406717980826105690264a26442, /* 2027 */
128'h0f230115c78300f10fa347090105c783, /* 2028 */
128'h02e78a63470d00e78e6301e1578300f1, /* 2029 */
128'hd06f6145b04505130000751770a27402, /* 2030 */
128'hd0efe42eadc5051300007517842a8b3f, /* 2031 */
128'hd8bff06f614570a265a2740285228a3f, /* 2032 */
128'h0113ebfff06f614505c170a241907402, /* 2033 */
128'h842a232130232291342322813823dc01, /* 2034 */
128'h22113c230028218006134581893284ae, /* 2035 */
128'he802c44a08282040061385a6e60ff0ef, /* 2036 */
128'h23813083f63ff0ef8522002cea2ff0ef, /* 2037 */
128'h24010113220139032281348323013403, /* 2038 */
128'h75974611cb8147a7d783000077978082, /* 2039 */
128'he40611418082cf3ff06f262585930000, /* 2040 */
128'ha70300e57763878e1041e703534000ef, /* 2041 */
128'h1007e78310a7a22310e1a02327051001, /* 2042 */
128'h4501808201418d5d91011782150260a2, /* 2043 */
128'hfc1ff0ef84aae426e822ec0611018082, /* 2044 */
128'h150202f407b33e800793470000ef842a, /* 2045 */
128'h610564a28d0502a7d533644260e29101, /* 2046 */
128'h00ef842af95ff0efe022e40611418082, /* 2047 */
128'h60a202f407b324078793000f47b74440, /* 2048 */
128'h1101808202a7d5330141910115026402, /* 2049 */
128'h892af63ff0ef84aae04ae426e822ec06, /* 2050 */
128'h24040413000f443702a48533412000ef, /* 2051 */
128'hfe856ee3f45ff0ef0405944a02855433, /* 2052 */
128'he426110180826105690264a2644260e2, /* 2053 */
128'h68048493842ae04aec06e822009894b7, /* 2054 */
128'hf0ef41240433854a89260084f3638922, /* 2055 */
128'h80826105690264a2644260e2f47dfa1f, /* 2056 */
128'h410007b7808200054503808200b50023, /* 2057 */
128'h4783410007378082020575130147c503, /* 2058 */
128'h07b7808200a70023dfe50207f7930147, /* 2059 */
128'h476d00e78623f8000713000782234100, /* 2060 */
128'h071300e78623470d0007822300e78023, /* 2061 */
128'h808200e788230200071300e78423fc70, /* 2062 */
128'h0146c7838082e31100054703410006b7, /* 2063 */
128'h2797b7e5050500e68023dfe50207f793, /* 2064 */
128'h97aa973e811100f5771334a787930000, /* 2065 */
128'h00f5802300e580a30007c78300074703, /* 2066 */
128'hf0efec068121842a002ce82211018082, /* 2067 */
128'hf0ef00914503f65ff0ef00814503fd1f, /* 2068 */
128'h00814503fb7ff0ef0ff47513002cf5df, /* 2069 */
128'h644260e2f43ff0ef00914503f4bff0ef, /* 2070 */
128'h892af406e84aec26f022717980826105, /* 2071 */
128'hf0ef0ff57513002c0089553b54e14461, /* 2072 */
128'h00914503f13ff0ef346100814503f81f, /* 2073 */
128'h694264e2740270a2fe9410e3f0bff0ef, /* 2074 */
128'h892af406e84aec26f022717980826145, /* 2075 */
128'h0ff57513002c0089553354e103800413, /* 2076 */
128'h4503ed1ff0ef346100814503f3fff0ef, /* 2077 */
128'h64e2740270a2fe9410e3ec9ff0ef0091, /* 2078 */
128'hf13ff0efec06002c1101808261456942, /* 2079 */
128'he9fff0ef00914503ea7ff0ef00814503, /* 2080 */
128'h842a4785e406e02211418082610560e2, /* 2081 */
128'h6797883dfefff0ef811135fd00b7d663, /* 2082 */
128'h60a2640200044503943e7da787930000, /* 2083 */
128'h439c3f27879300007797e69ff06f0141, /* 2084 */
128'h842e892aec4efc06f04af426f8227139, /* 2085 */
128'hb0ef19a505130000751702b7856384b2, /* 2086 */
128'h70e23ca7a32300007797c10d2501f0af, /* 2087 */
128'h771757fd8082612169e2790274a27442, /* 2088 */
128'h0000751785ca862600743af725230000, /* 2089 */
128'h00007797c50d2501fe5fa0ef16450513, /* 2090 */
128'h0000651785a604967563463238a7a823, /* 2091 */
128'h2923000077174785cdcfd0ef76450513, /* 2092 */
128'h099b00c4591bdd5ff0ef4521b77536f7, /* 2093 */
128'h993e0039791375e78793000067970009, /* 2094 */
128'hbf5d127010ef854edb7ff0ef00094503, /* 2095 */
128'he0221141bf953287ab23000077979c25, /* 2096 */
128'hd0efe4067345051300006517842a85aa, /* 2097 */
128'h8322f14025730ff0000f0000100fc82f, /* 2098 */
128'h830201410cc585930000559760a26402, /* 2099 */
128'h00007517404585930000659746051141, /* 2100 */
128'hc9112501d49fa0efe022e4062f450513, /* 2101 */
128'hd06f014160a264027185051300006517, /* 2102 */
128'h4605c26fd0ef7265051300006517c32f, /* 2103 */
128'h07850513000075177385859300006597, /* 2104 */
128'h7305051300006517c5112501d6bfa0ef, /* 2105 */
128'h0517bf6fd0ef5965051300006517b7e1, /* 2106 */
128'h77972807a32300007797e98505130000, /* 2107 */
128'h00054863842a8d0f90ef2607ad230000, /* 2108 */
128'h408005b3cf81439c26c7879300007797, /* 2109 */
128'hd06f014156c505130000651760a26402, /* 2110 */
128'h2501b6afb0ef00e5051300007517bb2f, /* 2111 */
128'h65974605bfb96de5051300006517c511, /* 2112 */
128'hc5112501c89fa0ef450133a585930000, /* 2113 */
128'hee1ff0ef8522b7816d85051300006517, /* 2114 */
128'hd39ff0efe40625011141900200000023, /* 2115 */
128'h80824501808224050513000f4537a001, /* 2116 */
128'h00756513157d631c1e07071300007717, /* 2117 */
128'h953e055e10d00513e308953600178693, /* 2118 */
128'he4328532ec06e822110102b506338082, /* 2119 */
128'h914ff0ef45816622c509842afd1ff0ef, /* 2120 */
128'h65171141808280826105644260e28522, /* 2121 */
128'h42000537af8fd0efe406672505130000, /* 2122 */
128'h8082450180820141450160a2eb5fc0ef, /* 2123 */
128'h808202f5553347a9b000257380824501, /* 2124 */
128'h05130000651785aa862e86b287361141, /* 2125 */
128'ha001c8bff0ef4505abcfd0efe40665e5, /* 2126 */
128'h07b3f57ff0efe406952e842ae0221141, /* 2127 */
128'h4505808201418d7d640260a295224080, /* 2128 */
128'hec26f022717980824505808245058082, /* 2129 */
128'h740270a20096186300c684bb842ef406, /* 2130 */
128'hc0efe432852285b280826145450164e2, /* 2131 */
128'h80824509bff92605200404136622e07f, /* 2132 */
128'h45018082808280828082450980824509, /* 2133 */
128'he822ec061101b8bff06f808245018082, /* 2134 */
128'h00d5043300d584b3003796934781e426, /* 2135 */
128'h80826105450164a2644260e200c79863, /* 2136 */
128'h65176090600c02e80363609800043803, /* 2137 */
128'h651785a286269fafd0ef5d2505130000, /* 2138 */
128'hbf5d0785a0019eafd0ef5ea505130000, /* 2139 */
128'he8a25ea5051300006517892ae0ca711d, /* 2140 */
128'he4a6ec86e862ec5ef05af456f852fc4e, /* 2141 */
128'h0a1300006a179bafd0ef44018b2ee466, /* 2142 */
128'h6c17fff949935deb8b9300006b975d6a, /* 2143 */
128'h0c9b996fd0ef85524ac15e2c0c130000, /* 2144 */
128'h9863448187ca98afd0ef855e85e60004, /* 2145 */
128'h974fd0ef856285e697cfd0ef85520364, /* 2146 */
128'h6517fd5417e3040502b49b63458187ca, /* 2147 */
128'h86b3a889450195afd0ef60a505130000, /* 2148 */
128'h40e9873300349713c689873e8a850084, /* 2149 */
128'h6390008586b3bf5d07a104856398e398, /* 2150 */
128'h0d6340e9873300359713c689873e8a85, /* 2151 */
128'h914fd0ef56c5051300006517058e02e6, /* 2152 */
128'h60e6557d908fd0ef5985051300006517, /* 2153 */
128'h6be27b027aa27a4279e2690664a66446, /* 2154 */
128'h7159bfa507a10585808261256ca26c42, /* 2155 */
128'he4ceeca6020005138aaa6a05fc56e0d2, /* 2156 */
128'he86aec66e8caf0a2f486f062f45ef85a, /* 2157 */
128'h0a134981b0fff0ef44818bb28b2ee46e, /* 2158 */
128'h8db300349793966c0c1300007c179c4a, /* 2159 */
128'h05130000651703749b6300fb0cb300fa, /* 2160 */
128'h6a0669a6694670a6740688efd0ef5665, /* 2161 */
128'h64e685da86266da26d426ce27c027ba2, /* 2162 */
128'hbadfe0efe33ff06f61657ae285567b42, /* 2163 */
128'he0ef892aba1fe0ef8d2aba7fe0ef842a, /* 2164 */
128'h6533010d1d1b0105151b0344f7b3b9bf, /* 2165 */
128'hb0238d4191011402150201a4643300a9, /* 2166 */
128'h0985a7dff0ef4521ef8100adb02300ac, /* 2167 */
128'h0485a6dff0ef0007c50397e20039f793, /* 2168 */
128'hf04af426f822fc06e032e42e7139b7ad, /* 2169 */
128'h892ab3ffe0ef842ab45fe0ef89aaec4e, /* 2170 */
128'h179b0105151bb33fe0ef84aab39fe0ef, /* 2171 */
128'h9101178265a2660215028fc18d450109, /* 2172 */
128'h9c63974e00e588330037971347818d5d, /* 2173 */
128'h863e69e2854e790274a270e2744200c7, /* 2174 */
128'h3703e3148ea907856314d79ff06f6121, /* 2175 */
128'he032e42e7139b7f100e830238f290008, /* 2176 */
128'hacdfe0ef89aaec4ef04af426f822fc06, /* 2177 */
128'he0ef84aaac1fe0ef892aac7fe0ef842a, /* 2178 */
128'h15028fc18d450109179b0105151babbf, /* 2179 */
128'h0037971347818d5d9101178265a26602, /* 2180 */
128'h74a270e2744200c79c63974e00e58833, /* 2181 */
128'h6314d01ff06f6121863e69e2854e7902, /* 2182 */
128'h00e830238f0900083703e3148e890785, /* 2183 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2184 */
128'h892aa4ffe0ef842aa55fe0ef89aaec4e, /* 2185 */
128'h179b0105151ba43fe0ef84aaa49fe0ef, /* 2186 */
128'h9101178265a2660215028fc18d450109, /* 2187 */
128'h9c63974e00e588330037971347818d5d, /* 2188 */
128'h863e69e2854e790274a270e2744200c7, /* 2189 */
128'he31402a686b307856314c89ff06f6121, /* 2190 */
128'h7139b7e100e8302302a7073300083703, /* 2191 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2192 */
128'h9cdfe0ef892a9d3fe0ef842a9d9fe0ef, /* 2193 */
128'h8d450109179b0105151b9c7fe0ef84aa, /* 2194 */
128'h47818d5d9101178265a2660215028fc1, /* 2195 */
128'h744200c79c63974e00e5883300379713, /* 2196 */
128'hf06f6121863e69e2854e790274a270e2, /* 2197 */
128'he31402a6d6b3078563144505e111c0df, /* 2198 */
128'h7139b7d100e8302302a7573300083703, /* 2199 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2200 */
128'h94dfe0ef892a953fe0ef842a959fe0ef, /* 2201 */
128'h8d450109179b0105151b947fe0ef84aa, /* 2202 */
128'h47818d5d9101178265a2660215028fc1, /* 2203 */
128'h744200c79c63974e00e5883300379713, /* 2204 */
128'hf06f6121863e69e2854e790274a270e2, /* 2205 */
128'h8f4900083703e3148ec907856314b8df, /* 2206 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2207 */
128'he0ef842a8e1fe0ef89aaec4ef04af426, /* 2208 */
128'h151b8cffe0ef84aa8d5fe0ef892a8dbf, /* 2209 */
128'h65a2660215028fc18d450109179b0105, /* 2210 */
128'h00e588330037971347818d5d91011782, /* 2211 */
128'h854e790274a270e2744200c79c63974e, /* 2212 */
128'h8ee907856314b15ff06f6121863e69e2, /* 2213 */
128'h7139b7f100e830238f6900083703e314, /* 2214 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2215 */
128'h85dfe0ef892a863fe0ef842a869fe0ef, /* 2216 */
128'h8cc90109179b0105151b857fe0ef84aa, /* 2217 */
128'h47018fc59081178265a2660214828fc1, /* 2218 */
128'h744200c71c6396ae00d9883300371693, /* 2219 */
128'hf06f6121863a69e2854e790274a270e2, /* 2220 */
128'hbfc9070500a83023e28800f70533a9df, /* 2221 */
128'hf0a20ca5051300006517892ae8ca7159, /* 2222 */
128'heca6f486f062f45ef85afc56e0d2e4ce, /* 2223 */
128'h00006a17c99fc0ef44018b3289aeec66, /* 2224 */
128'h00006c170bcb8b9300006b970b4a0a13, /* 2225 */
128'h4493c77fc0ef855204000a930c4c0c13, /* 2226 */
128'h40900cb3c69fc0ef8885855e85a2fff4, /* 2227 */
128'h186397ce00f905b30036179314fd4601, /* 2228 */
128'hc0ef856285a2c4bfc0efe43285520566, /* 2229 */
128'he12984aaa03ff0ef854a85ce6622c43f, /* 2230 */
128'hc0ef0d25051300006517fb541be32405, /* 2231 */
128'h6a0669a664e669468526740670a6c23f, /* 2232 */
128'h7693808261656ce27c027ba27b427ae2, /* 2233 */
128'hbf590605e198e3988726c29187660016, /* 2234 */
128'h05130000651784aaeca67159bfc154fd, /* 2235 */
128'hf45ef85afc56e0d2e4cee8caf0a2ff65, /* 2236 */
128'hc0ef44018ab2892ee86af486ec66f062, /* 2237 */
128'h0b1300006b17fde9899300006997bc3f, /* 2238 */
128'h0c1300006c17326b8b9300006b97326b, /* 2239 */
128'h854e04000a13fdec8c9300006c97fd6c, /* 2240 */
128'h85a2000bbd03cba500147793b91fc0ef, /* 2241 */
128'h00361793fffd45134601b7ffc0ef8562, /* 2242 */
128'hc0efe432854e05561c6397ca00f485b3, /* 2243 */
128'h852685ca6622b5bfc0ef856685a2b63f, /* 2244 */
128'h6517fb441ae32405e5298d2a91bff0ef, /* 2245 */
128'h856a740670a6b3bfc0effea505130000, /* 2246 */
128'h7c027ba27b427ae26a0669a6694664e6, /* 2247 */
128'h7693bf49000b3d03808261656d426ce2, /* 2248 */
128'hb7790605e198e398872ac291876a0016, /* 2249 */
128'h051300006517842ae8a2711db7e15d7d, /* 2250 */
128'he862ec5ef05af456f852e0cae4a6f065, /* 2251 */
128'h6917ad7fc0ef4c018ab284aefc4eec86, /* 2252 */
128'h6b97efab0b1300006b17ef2909130000, /* 2253 */
128'hab5fc0ef854a10000a13f02b8b930000, /* 2254 */
128'h008c1713aa9fc0ef855a85ce000c099b, /* 2255 */
128'h8fd9018c17130187e7b38fd9010c1793, /* 2256 */
128'h030c17138fd9028c17138fd9020c1713, /* 2257 */
128'h06b30036171346018fd9038c17138fd9, /* 2258 */
128'ha65fc0efe432854a05561763972600e4, /* 2259 */
128'hf0ef852285a66622a5dfc0ef855e85ce, /* 2260 */
128'h00006517f94c19e30c05e91d89aa81df, /* 2261 */
128'h64a6854e644660e6a3dfc0efeec50513, /* 2262 */
128'h61256c426be27b027aa27a4279e26906, /* 2263 */
128'h7119bff159fdb74d0605e29ce31c8082, /* 2264 */
128'hf0caf8a2e1c505130000651784aaf4a6, /* 2265 */
128'hf06af466f862fc5ee0dae4d6e8d2ecce, /* 2266 */
128'h6a179e7fc0ef44018b32892eec6efc86, /* 2267 */
128'h0b93e0ac8c9300006c97e02a0a130000, /* 2268 */
128'he08d0d1300006d1703f00c13498507f0, /* 2269 */
128'hc0ef856685a29bbfc0ef855208000a93, /* 2270 */
128'h4601008995b300e99733408b873b9b3f, /* 2271 */
128'h855205661a6397ca00f486b300361793, /* 2272 */
128'h6622987fc0ef856a85a298ffc0efe432, /* 2273 */
128'h1be32405e1398daaf46ff0ef852685ca, /* 2274 */
128'h70e6967fc0efe165051300006517fb54, /* 2275 */
128'h6b066aa66a4669e6790674a6856e7446, /* 2276 */
128'h6663808261096de27d027ca27c427be2, /* 2277 */
128'hbfe5e298e398bf610605e28ce38c008c, /* 2278 */
128'h05130000651784aaf4a67119b7f15dfd, /* 2279 */
128'hfc5ee0dae4d6e8d2eccef0caf8a2d365, /* 2280 */
128'h44018b32892eec6efc86f06af466f862, /* 2281 */
128'h00006c97d1ca0a1300006a17901fc0ef, /* 2282 */
128'h6d1703f00c13498507f00b93d24c8c93, /* 2283 */
128'h8d5fc0ef855208000a93d22d0d130000, /* 2284 */
128'h00f997b3408b87bb8cdfc0ef856685a2, /* 2285 */
128'h17134601fff6c693fff7c793008996b3, /* 2286 */
128'he432855205661a63974a00e485b30036, /* 2287 */
128'h85ca6622899fc0ef856a85a28a1fc0ef, /* 2288 */
128'hfb5417e32405e1398daae58ff0ef8526, /* 2289 */
128'h744670e6879fc0efd285051300006517, /* 2290 */
128'h7be26b066aa66a4669e6790674a6856e, /* 2291 */
128'h008c6663808261096de27d027ca27c42, /* 2292 */
128'h5dfdbfe5e19ce31cbf610605e194e314, /* 2293 */
128'hc48505130000651784aaf4a67119b7f1, /* 2294 */
128'hf862fc5ee0dae4d6e8d2eccef0caf8a2, /* 2295 */
128'hc0ef44018a32892eec6efc86f06af466, /* 2296 */
128'h0c1300006c17c2e9899300006997813f, /* 2297 */
128'h03f00b9308100b134d0507f00a93c36c, /* 2298 */
128'h85a2fe6fc0ef854ec30c8c9300006c97, /* 2299 */
128'h17b3408b07bb408a873bfdefc0ef8562, /* 2300 */
128'h00fd17b30024079b8f5d00ed173300fd, /* 2301 */
128'h4601fff7c313fff748938fd5008d16b3, /* 2302 */
128'h854e05461c6396ca00d4853300361693, /* 2303 */
128'h6622f96fc0ef856685a2f9efc0efe432, /* 2304 */
128'h07932405ed298daad56ff0ef852685ca, /* 2305 */
128'hc0efc225051300006517f8f41be30800, /* 2306 */
128'h6a4669e6790674a6856e744670e6f72f, /* 2307 */
128'h61096de27d027ca27c427be26b066aa6, /* 2308 */
128'h00081363859a008bea63001678138082, /* 2309 */
128'hfe081be385c6b7610605e10ce28c85be, /* 2310 */
128'h6517892af0ca7119bf755dfdbfc585ba, /* 2311 */
128'hf06af466fc5ee8d2ecceb32505130000, /* 2312 */
128'h89aef862e0dae4d6f4a6f8a2fc86ec6e, /* 2313 */
128'hb18a0a1300006a17efcfc0ef4b81e032, /* 2314 */
128'hb28d0d1300006d17b20c8c9300006c97, /* 2315 */
128'h85524401003b949b01779c3347854da1, /* 2316 */
128'hec4fc0ef856685da00848b3bed0fc0ef, /* 2317 */
128'h00e908330036171367824601fffc4a93, /* 2318 */
128'h85daea6fc0efe432855206f61063974e, /* 2319 */
128'hc5eff0ef854a85ce6622e9efc0ef856a, /* 2320 */
128'h07932b85fbb41be38c562405e9318b2a, /* 2321 */
128'hc0efb225051300006517fafb90e30400, /* 2322 */
128'h6a4669e6790674a6855a744670e6e72f, /* 2323 */
128'h61096de27d027ca27c427be26b066aa6, /* 2324 */
128'h3023e30c85d6e11185e2001675138082, /* 2325 */
128'hf8cafca67175b7e95b7db749060500b8, /* 2326 */
128'hecd6f0d2698502000513892e84aaf4ce, /* 2327 */
128'hf46ef86ae122e506fc66e0e2e4dee8da, /* 2328 */
128'h0c1300006c174a01862ff0ef4a81e032, /* 2329 */
128'h8b26eb2c8c9300006c979c4989936f6c, /* 2330 */
128'h956396da003d969367824d214d818bca, /* 2331 */
128'hed45842aba2ff0ef852685ca866e04fd, /* 2332 */
128'hdc4fc0efa9c5051300006517020a0863, /* 2333 */
128'h6ae67a0679a6794674e6640a60aa8522, /* 2334 */
128'h808261497da27d427ce26c066ba66b46, /* 2335 */
128'h842a8defe0efec36b7758ba68b4a4a05, /* 2336 */
128'h8ccfe0efe42a8d2fe0efe82a8d8fe0ef, /* 2337 */
128'h8c510106161b8d5d0105151b664267a2, /* 2338 */
128'hbb23000067978d4166e2910114021502, /* 2339 */
128'h86330006c683018786b34781e28864a7, /* 2340 */
128'hffa795e300d600230ff6f693078500fb, /* 2341 */
128'h879bf8dfe0ef4521ef910ba1033df7b3, /* 2342 */
128'he0ef0007c50397e68b8d00078a9b001a, /* 2343 */
128'hf4cef8ca7175bfa1547dbf0d0d85f79f, /* 2344 */
128'hecd6fca66a050200051389ae892af0d2, /* 2345 */
128'hf46ee122e506f86afc66e0e2e4dee8da, /* 2346 */
128'h8493000064974a81f43fe0ef4b018cb2, /* 2347 */
128'h8bcad92d0d1300006d179c4a0a135de4, /* 2348 */
128'h956397de00fc06b3003d97934d818c4e, /* 2349 */
128'he579842aa82ff0ef854a85ce866e059d, /* 2350 */
128'hca4fc0ef97c5051300006517020a8863, /* 2351 */
128'h6ae67a0679a6794674e6640a60aa8522, /* 2352 */
128'h808261497da27d427ce26c066ba66b46, /* 2353 */
128'hfbdfd0efe836ec3eb7758c4a8bce4a85, /* 2354 */
128'hd0efe02afb1fd0efe42afb7fd0ef842a, /* 2355 */
128'h8d590106161b0105151b67026622fabf, /* 2356 */
128'hbf23000067978d419101140215028c51, /* 2357 */
128'h93c117c20004d783e38866c267e252a7, /* 2358 */
128'h00f6912393c117c20024d78300f69023, /* 2359 */
128'h0064d78300f6922393c117c20044d783, /* 2360 */
128'h4521ef91034df7b300f6932393c117c2, /* 2361 */
128'h97ea8b8d00078b1b001b079be57fe0ef, /* 2362 */
128'hb789547dbf290d85e43fe0ef0007c503, /* 2363 */
128'he122fff586138932f8ca717580826505, /* 2364 */
128'h05130000651785aa962a84ae842afca6, /* 2365 */
128'hfc66e0e2e4dee8daecd6f0d2f4ce89e5, /* 2366 */
128'h0044d793ba8fc0efec36e506f46ef86a, /* 2367 */
128'h4a81e43e99a20034d793e83e0014d993, /* 2368 */
128'h8b9300006b97886b0b1300006b174485, /* 2369 */
128'h8c9300006c97886c0c1300006c17886b, /* 2370 */
128'h8d9300006d9788ed0d1300006d17886c, /* 2371 */
128'h651702997863436a0a1300006a1788ed, /* 2372 */
128'h8556640a60aab4afc0ef882505130000, /* 2373 */
128'h6c066ba66b466ae67a0679a6794674e6, /* 2374 */
128'hc0ef855a85a6808261497da27d427ce2, /* 2375 */
128'h8562b16fc0ef855e85ca00090663b22f, /* 2376 */
128'h852265a2b08fc0ef856a85e6b10fc0ef, /* 2377 */
128'h010a2783af8fc0ef856eed15920ff0ef, /* 2378 */
128'h00006517c58d000a358302f749636762, /* 2379 */
128'h85ce6642008a3783adcfc0ef80450513, /* 2380 */
128'hac4fc0ef7f4505130000551797828522, /* 2381 */
128'hab4fc0ef5ac5051300005517b7e94a89, /* 2382 */
128'h7e05051300005517c62a7139bfa10485, /* 2383 */
128'h0597be7fe0efec4ef04af426f822fc06, /* 2384 */
128'hc0ef7da5051300005517fe6585930000, /* 2385 */
128'ha74fc0ef7e45051300005517006ca82f, /* 2386 */
128'ha64fc0ef7e4505130000551704000593, /* 2387 */
128'h00006517a58fc0ef8005051300006517, /* 2388 */
128'h5385051300005517a4cfc0ef82450513, /* 2389 */
128'h95b3497901f499934441a3efc0ef4485, /* 2390 */
128'he49ff0ef240501358533460546850084, /* 2391 */
128'h612169e2790274a2744270e2ff2417e3, /* 2392 */
128'h46814881470100c5131b460580828082, /* 2393 */
128'h000780234000081387f245a901f61e13, /* 2394 */
128'h802397aa0007802397aa0007802397aa, /* 2395 */
128'h02b71d632705fe0813e397aa387d0007, /* 2396 */
128'h86b33e800513c00026f38e15c0202673, /* 2397 */
128'h45bb02c747334000059302a687334116, /* 2398 */
128'h05130000551702a7473302a767b302b3, /* 2399 */
128'h28f3c02026f3fac710e399efc06f7be5, /* 2400 */
128'h4505f7bff0ef4501e4061141bf51c000, /* 2401 */
128'hf69ff0ef4511f6fff0ef4509f75ff0ef, /* 2402 */
128'h6697bff1f5dff0ef4541f63ff0ef4521, /* 2403 */
128'h6a630ae50963429c4729262686930000, /* 2404 */
128'h871bc30507f7f7130ce51b63472108a7, /* 2405 */
128'h0706450387b722e62f2300006617fff7, /* 2406 */
128'h6785429800e79023f207071b776597ba, /* 2407 */
128'h2b2300006617c007071b670504f74863, /* 2408 */
128'h87938007071376654503a737650520e6, /* 2409 */
128'h55830af84363f206061bf7f50813c007, /* 2410 */
128'h96e30709278500b7102391c115c21007, /* 2411 */
128'h1cf72c2300006717f807879b6785fea7, /* 2412 */
128'hef1c879deb1407f7f6934503c737429c, /* 2413 */
128'hf793b7a507f0071300e5056347358082, /* 2414 */
128'he5137665b7491af7272300006717f807, /* 2415 */
128'hf206061b450388b745810017971307f7, /* 2416 */
128'h10239746b78dfde900f5546300270813, /* 2417 */
128'h66170017871bb7e587424585278500c7, /* 2418 */
128'h670597ba45038737078616e629230000, /* 2419 */
128'hb73d00a79023914115428d59f0070713, /* 2420 */
128'hc007879b6785955fe06fb79d00c71023, /* 2421 */
128'he4064503c7b7114114f7202300006717, /* 2422 */
128'h6705ef98020007130007b823e7984729, /* 2423 */
128'h83370713f79481470693f39480070693, /* 2424 */
128'h4741e3b831300713ff9830000713fb98, /* 2425 */
128'h0713f7b818000713f3b831000713efb8, /* 2426 */
128'h02800713e3d8472dffb84715fbb87800, /* 2427 */
128'h373710e7b02372d7071300202737ebd8, /* 2428 */
128'h071300e9373710e7b42354f7071300e0, /* 2429 */
128'hbc236e87071300e1e73710e7b82374f7, /* 2430 */
128'hb4230aa7071312e7b02300aa073710e7, /* 2431 */
128'hb73712e7b8235007071300aa573712e7, /* 2432 */
128'h06930055573712e7bc23aaa7071300aa, /* 2433 */
128'h073714e7b4235ff7071314d7b0235557, /* 2434 */
128'h14e7bc23177d14d7b823f55706930056, /* 2435 */
128'h5ff7071316d7b0235557069300ff5737, /* 2436 */
128'h16d7b823f55706930100073716e7b423, /* 2437 */
128'h06130000161716e7bc234503e5b7177d, /* 2438 */
128'h8e334701489100c5881345314781c266, /* 2439 */
128'h070500ee03330006c68300e606b300b7, /* 2440 */
128'h4701fea714e300d3002307e6f6938285, /* 2441 */
128'h1be307050006802300e306b301078333, /* 2442 */
128'h4503f7b7f36906318007871307c1ff17, /* 2443 */
128'h070500d700238107879356fd80078713, /* 2444 */
128'h0007b02345070737450407b7fef71de3, /* 2445 */
128'he39875e147094503c7b7fee79de307a1, /* 2446 */
128'h0e9306b0089308058593786145038637, /* 2447 */
128'h07bb4503ae370800031308000f130750, /* 2448 */
128'h8fcd0807e5134107d79b0107979b0106, /* 2449 */
128'h02e8c763470186b293c1914117c21542, /* 2450 */
128'h10060613fe671ae30689270500f69023, /* 2451 */
128'hc7b760a20ee000ef02800513fdc617e3, /* 2452 */
128'h902300eec56380820141e39847054503, /* 2453 */
128'he02211418082b7f100a69023bfc901e6, /* 2454 */
128'h014160a264028522f36fe0ef842ae406, /* 2455 */
128'h00044503842ae406e0221141cbfff06f, /* 2456 */
128'hfd1ff0ef040580820141640260a2e509, /* 2457 */
128'h079b440184aaf406ec26f0227179b7f5, /* 2458 */
128'h8082614564e2740270a200b7c7630004, /* 2459 */
128'hfa1ff0ef0405e42e0007c503008487b3, /* 2460 */
128'h80820ff0051380820ff00513bff165a2, /* 2461 */
128'h7513842ae022715d8082808280824501, /* 2462 */
128'he0c2fc3ef83af436f032ec2ee4060ff5, /* 2463 */
128'h80826161640260a28522f6bff0efe4c6, /* 2464 */
128'h4529e90900044503842ae406e0221141, /* 2465 */
128'h0405808201414501640260a2f4dff0ef, /* 2466 */
128'h4f878793000057971101b7d5f3dff0ef, /* 2467 */
128'h189be44ae826ec220007b30300034e37, /* 2468 */
128'h478146014e8103658593000015970045, /* 2469 */
128'hc8039ffe0e131ff00f9362994f3d4681, /* 2470 */
128'h0003841b0188181b07f8739305850005, /* 2471 */
128'h0029149b00f7f9130005c7034188581b, /* 2472 */
128'hfb6301e91e6302a684b38e5900971733, /* 2473 */
128'h070e97268311ff1787130054f9630117, /* 2474 */
128'h00f7e79300fff86307854601e310971a, /* 2475 */
128'h347d058500084363478106850317ee63, /* 2476 */
128'h53639eba070593011702fff3871bf855, /* 2477 */
128'hfd63661902a687b3f9de75e305850008, /* 2478 */
128'h00f7f713a01d4681971a0037971302c7, /* 2479 */
128'h971a070e97268311ff17871301e71a63, /* 2480 */
128'h0721068500073023b76d07854601e310, /* 2481 */
128'h4107879300005797b7e197aafea69ce3, /* 2482 */
128'hb02300e036b772d7071300202737639c, /* 2483 */
128'h071310d7b42300e9373754f6869310e7, /* 2484 */
128'h646212e7b02310d7bc2310e7b82374f7, /* 2485 */
128'h692264c212e7b4236e87071300e1e737, /* 2486 */
128'h1582892e02100793f84a715d80826105, /* 2487 */
128'hec56920195be160289b29181f44e07ea, /* 2488 */
128'h8aaae062e45ee85af052fc26e0a2e486, /* 2489 */
128'h74e2640660a606f962636785a53fd0ef, /* 2490 */
128'h61616c026ba26b426ae27a0279a27942, /* 2491 */
128'he4afe0ef910145a115020089053b8082, /* 2492 */
128'h4481bc7fb0ef020c5c13855202041c13, /* 2493 */
128'he0ef048545890007c50397d6009c07b3, /* 2494 */
128'hb0ef855eff6494e3badfb0ef8552e28f, /* 2495 */
128'h00004a174401b74dfb346fe32441ba3f, /* 2496 */
128'hb7dde7ab8b9300005b974b412d4a0a13, /* 2497 */
128'h440007b78082e388440007b791011502, /* 2498 */
128'h6b880007b823440007b7808225016388, /* 2499 */
128'hf7b7808225017b88440007b780822501, /* 2500 */
128'h959b8ed192518efd165200c6969b00ff, /* 2501 */
128'h8ecd8dfd0185159b7f0007b78ecd01f5, /* 2502 */
128'h4400063747812501f7942681440007b7, /* 2503 */
128'h440006b73e80079300a6ef630007869b, /* 2504 */
128'h7388440007b7ffe537fdc3198b097a98, /* 2505 */
128'hf61407850006e68396ba002796938082, /* 2506 */
128'hfc26e0a20210091347cdf84a715dbfc1, /* 2507 */
128'h44814401c43ee486e85aec56f052f44e, /* 2508 */
128'h07bb1ff009935b61096a5afd00b00a37, /* 2509 */
128'h4509458102700613041006930038009a, /* 2510 */
128'h07938726240503551f63f5dff0efc63e, /* 2511 */
128'h802396ca00f556339281020716930380, /* 2512 */
128'hfc89f1e324a1ff6796e3270537e100c6, /* 2513 */
128'h6b426ae27a0279a2794274e2640660a6, /* 2514 */
128'h0513000055171141b7d9440180826161, /* 2515 */
128'h00005517f6bff0efa5dfb0efe4060c65, /* 2516 */
128'he1c5051300000517a4dfb0ef0d450513, /* 2517 */
128'h551740a005b360a200055c63f36f70ef, /* 2518 */
128'h014160a2a29fb06f0141be2505130000, /* 2519 */
128'hb64fe06f1545051300005517d8cfe06f, /* 2520 */
128'he456e852ec4ef04af426f822fc067139, /* 2521 */
128'he0ef0925051300005517b1cfe0efe05a, /* 2522 */
128'h00005917440009b79a7ff0ef4401b42f, /* 2523 */
128'h059b639097ce00341793449508c90913, /* 2524 */
128'h70effe9416e39cbfb0ef0405854a0004, /* 2525 */
128'h440004b7174b0b1300005b174901f9ff, /* 2526 */
128'h078a0a1300005a17068a8a9300005a97, /* 2527 */
128'he09c090585560007c783016907b34991, /* 2528 */
128'hb823987fb0ef8622240125816080608c, /* 2529 */
128'hfd391be3979fb0ef25818552688c0004, /* 2530 */
128'h371702f7646347190054579b0ff47413, /* 2531 */
128'h878297ba439c97ba078a59a707130000, /* 2532 */
128'he0ef8522949fb0ef0385051300005517, /* 2533 */
128'h935fb0ef0345051300005517a001ce2f, /* 2534 */
128'h0305051300005517b7f5ec7ff0ef8522, /* 2535 */
128'h00005517bfe1e6eff0ef8522921fb0ef, /* 2536 */
128'h5517b7d981cf80ef90dfb0ef02c50513, /* 2537 */
128'hbf55f6aff0ef8fbfb0ef02a505130000, /* 2538 */
128'h00000000000000000000000000000000, /* 2539 */
128'h00000000000000000000000000000000, /* 2540 */
128'h00000000000000000000000000000000, /* 2541 */
128'h00000000000000000000000000000000, /* 2542 */
128'h00000000000000000000000000000000, /* 2543 */
128'h08082828282828080808080808080808, /* 2544 */
128'h08080808080808080808080808080808, /* 2545 */
128'h101010101010101010101010101010a0, /* 2546 */
128'h10101010101004040404040404040404, /* 2547 */
128'h01010101010101010141414141414110, /* 2548 */
128'h10101010100101010101010101010101, /* 2549 */
128'h02020202020202020242424242424210, /* 2550 */
128'h08101010100202020202020202020202, /* 2551 */
128'h00000000000000000000000000000000, /* 2552 */
128'h00000000000000000000000000000000, /* 2553 */
128'h101010101010101010101010101010a0, /* 2554 */
128'h10101010101010101010101010101010, /* 2555 */
128'h01010101010101010101010101010101, /* 2556 */
128'h02010101010101011001010101010101, /* 2557 */
128'h02020202020202020202020202020202, /* 2558 */
128'h02020202020202021002020202020202, /* 2559 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2560 */
128'hfd469501a83046134787c62af57c0faf, /* 2561 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2562 */
128'h49b40821a679438efd9871936b901122, /* 2563 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2564 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2565 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2566 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2567 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2568 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2569 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2570 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2571 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2572 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2573 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2574 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2575 */
128'h0c07020d08030e09040f0a05000b0601, /* 2576 */
128'h020f0c090603000d0a0704010e0b0805, /* 2577 */
128'h09020b040d060f08010a030c050e0700, /* 2578 */
128'h6c5f7465735f64735f63736972776f6c, /* 2579 */
128'h6e67696c615f64730000000000006465, /* 2580 */
128'h645f6b6c635f64730000000000000000, /* 2581 */
128'h69747465735f64730000000000007669, /* 2582 */
128'h735f646d635f6473000000000000676e, /* 2583 */
128'h74657365725f64730000000074726174, /* 2584 */
128'h6e636b6c625f64730000000000000000, /* 2585 */
128'h69736b6c625f64730000000000000074, /* 2586 */
128'h6f656d69745f6473000000000000657a, /* 2587 */
128'h655f7172695f64730000000000007475, /* 2588 */
128'h5f63736972776f6c000000000000006e, /* 2589 */
128'h00000000646d635f74726174735f6473, /* 2590 */
128'h746e695f746961775f63736972776f6c, /* 2591 */
128'h000000000067616c665f747075727265, /* 2592 */
128'h00007172695f64735f63736972776f6c, /* 2593 */
128'h695f646d635f64735f63736972776f6c, /* 2594 */
128'h5f63736972776f6c0000000000007172, /* 2595 */
128'h007172695f646e655f617461645f6473, /* 2596 */
128'h0000000087fea2880000000087fee4a0, /* 2597 */
128'h004c4b40004c4b400030000020000000, /* 2598 */
128'h6d6d5f6472616f62000000020000ffff, /* 2599 */
128'h0000000087fe4ea40064637465675f63, /* 2600 */
128'h0000000087fe4d100000000087fe4ab2, /* 2601 */
128'h00000000000000000000000000000000, /* 2602 */
128'hffffb586ffffb582ffffb582ffffb55c, /* 2603 */
128'hffffb58affffb58affffb58affffb58a, /* 2604 */
128'h0000000087fee7c80000000087fee7b8, /* 2605 */
128'h0000000087fee7f00000000087fee7d8, /* 2606 */
128'h0000000087fee8200000000087fee808, /* 2607 */
128'h0000000087fee8500000000087fee838, /* 2608 */
128'h0000000087fee8800000000087fee868, /* 2609 */
128'h0000000087fee8b00000000087fee898, /* 2610 */
128'h40040300400402004004010040040000, /* 2611 */
128'h40050000400405004004040140040400, /* 2612 */
128'h30000000000000030000000040050100, /* 2613 */
128'h60000000000000053000000000000001, /* 2614 */
128'h70000000000000027000000000000004, /* 2615 */
128'h00000001400000007000000000000000, /* 2616 */
128'h00000005000000012000000000000006, /* 2617 */
128'h20000000000000020000000040000000, /* 2618 */
128'h00000000100000000000000100000000, /* 2619 */
128'h1e19140f0d0c0a000000000000000000, /* 2620 */
128'h000186a00000271050463c37322d2823, /* 2621 */
128'h017d7840017d784000989680000f4240, /* 2622 */
128'h031975000319750002faf080018cba80, /* 2623 */
128'h02faf08005f5e10002faf080017d7840, /* 2624 */
128'h00000020000000000bebc2000c65d400, /* 2625 */
128'h00000200000001000000008000000040, /* 2626 */
128'h00002000000010000000080000000400, /* 2627 */
128'h0000c000000080000000600000004000, /* 2628 */
128'h37363534333231300002000000010000, /* 2629 */
128'h2043534952776f4c4645444342413938, /* 2630 */
128'h746f6f622d7520646573696d696e696d, /* 2631 */
128'h00000000647261432d445320726f6620, /* 2632 */
128'h18100000000000002060fcfc60200000, /* 2633 */
128'h30303030fc783000000000001018fcfc, /* 2634 */
128'h00003078fc3030303030300000003030, /* 2635 */
128'hb2847800000078848282828282847800, /* 2636 */
128'h828282828282fe0000007884b2fafafa, /* 2637 */
128'h0000fe86cefab2face86fe000000fe82, /* 2638 */
128'h700000000080c0e0f0f8fcf8f0e0c080, /* 2639 */
128'h181e0600000000000000000070f8f8f8, /* 2640 */
128'h3030303060e080000000000030303030, /* 2641 */
128'h303030300000000000061e1830303030, /* 2642 */
128'h00fefe0000000000000000000080e060, /* 2643 */
128'h30303030303030303030303000000000, /* 2644 */
128'h303030303030303030fefe0000000000, /* 2645 */
128'h303e3e30303030300000000000fefe30, /* 2646 */
128'h3030303030f0f0303030303030303030, /* 2647 */
128'h00fefe003030303030fefe3030303030, /* 2648 */
128'h66b298cc66b298cc00fefe0000fefe00, /* 2649 */
128'hcccccccccccccccccccccccc66b298cc, /* 2650 */
128'he0e0e0e0aad4aad4aad4aad4aad4aad4, /* 2651 */
128'h1e1ee0e0e0e0e0e0fefefefefefee0e0, /* 2652 */
128'he0e0e0e0e0e0e0e0e0e0e0e01e1e1e1e, /* 2653 */
128'h00000000000000000000e0e0e0e0e0e0, /* 2654 */
128'h1e1e000000000000fefefefefefe0000, /* 2655 */
128'he0e0e0e0e0e00000000000001e1e1e1e, /* 2656 */
128'h20200000000000000000000000000000, /* 2657 */
128'h00000000505028000000200020202020, /* 2658 */
128'h00005050fc5028fc2828000000000000, /* 2659 */
128'ha84800000020f0a8283060a0a8782000, /* 2660 */
128'ha8a878505020000000004854342850b0, /* 2661 */
128'h00000000000000008040400000006c90, /* 2662 */
128'h10204000000408101010101010080400, /* 2663 */
128'ha87070a8200000000040201010101010, /* 2664 */
128'h000000202020f8202020000000000020, /* 2665 */
128'h00000000804040000000000000000000, /* 2666 */
128'h0000000000000000000000000000f800, /* 2667 */
128'h00804040402020101010080000004000, /* 2668 */
128'h60200000000070888888888888700000, /* 2669 */
128'h40201088887000000000702020202020, /* 2670 */
128'h0000708808083008887000000000f880, /* 2671 */
128'h80f80000000018107890505030100000, /* 2672 */
128'h8888f08090700000000070880808f080, /* 2673 */
128'h000020202020201090f8000000007088, /* 2674 */
128'h88700000000070888888708888700000, /* 2675 */
128'h00000020000000000000704808788888, /* 2676 */
128'h00202000000020000000000000002000, /* 2677 */
128'h00000000000004081020402010080400, /* 2678 */
128'h100804081020400000000000f80000f8, /* 2679 */
128'h00002000202010888870000000004020, /* 2680 */
128'h2020000000007880b8a8a89888700000, /* 2681 */
128'h4848704848f000000000cc4878505030, /* 2682 */
128'h0000708880808080887800000000f048, /* 2683 */
128'h48f800000000f0484848484848f00000, /* 2684 */
128'h4050705048f800000000f84840507050, /* 2685 */
128'h00003048889c8080483800000000e040, /* 2686 */
128'h20f800000000cc484848784848cc0000, /* 2687 */
128'h10101010107c00000000f82020202020, /* 2688 */
128'h0000ec485050605048ec000000e09010, /* 2689 */
128'hd8d800000000fc444040404040e00000, /* 2690 */
128'h5858686848dc00000000a8a8a8a8d8d8, /* 2691 */
128'h0000708888888888887000000000e848, /* 2692 */
128'h887000000000e0404040704848f00000, /* 2693 */
128'h4850704848f0000000187098e8888888, /* 2694 */
128'h0000f08808106080887800000000ec48, /* 2695 */
128'h48cc00000000702020202020a8f80000, /* 2696 */
128'h3050504848cc00000000304848484848, /* 2697 */
128'h00005050505070a8a8a8000000002020, /* 2698 */
128'h50d800000000d8505020205050d80000, /* 2699 */
128'h4020201090f800000000702020202050, /* 2700 */
128'h0038202020202020202038000000f848, /* 2701 */
128'h10107000000008101010202040404000, /* 2702 */
128'h00000000005020000070101010101010, /* 2703 */
128'hfc000000000000000000000000000000, /* 2704 */
128'h00000000000000000000000000002000, /* 2705 */
128'h4848704040c0000000003c4838483000, /* 2706 */
128'h00003840404838000000000000007048, /* 2707 */
128'h0000000000003c484848380808180000, /* 2708 */
128'h20207820201c00000000384078483000, /* 2709 */
128'h3844784030483c000000000000007820, /* 2710 */
128'h002000000000ec484848704040c00000, /* 2711 */
128'h10103000001000000000702020206000, /* 2712 */
128'h0000ec4870505c4040c00000e0101010, /* 2713 */
128'h000000000000f8202020202020e00000, /* 2714 */
128'h4848f000000000000000a8a8a8a8f000, /* 2715 */
128'h0000304848483000000000000000ec48, /* 2716 */
128'h00000000e04070484848f00000000000, /* 2717 */
128'h4060d800000000001c08384848483800, /* 2718 */
128'h0000780830407800000000000000e040, /* 2719 */
128'h00000000000018202020702020000000, /* 2720 */
128'h5048ec000000000000003c484848d800, /* 2721 */
128'h0000505070a8a8000000000000002030, /* 2722 */
128'h000000000000d8502050d80000000000, /* 2723 */
128'h2010780000000000c02020305048ec00, /* 2724 */
128'h00181010101020101010180000007820, /* 2725 */
128'h20206000101010101010101010101010, /* 2726 */
128'h000000000018a4400060202020201020, /* 2727 */
128'h00ff018d00fa00ff0000000000000000, /* 2728 */
128'h00d600ff00ff00ff01a600e900ff00ff, /* 2729 */
128'h00ff00ff00ff0182028201ab02820183, /* 2730 */
128'h00ff00ff0182028201b10282018300cc, /* 2731 */
128'h00ff0184020101bc0201018300c400ff, /* 2732 */
128'h00ff03020201c802010200ba00ff00ff, /* 2733 */
128'h0182020101cb0282010100b500ff00ff, /* 2734 */
128'h020101d20201018200ae00ff00ff00ff, /* 2735 */
128'h01d50201018200aa00ff00ff00ff0182, /* 2736 */
128'h00ff01e100a500ff00ff00ff01820201, /* 2737 */
128'hff00ff00ff03020201e5009f00ff00ff, /* 2738 */
128'hff00ff00ff03020201e6020102009a00, /* 2739 */
128'h00ff00ff03020201eb02010182009600, /* 2740 */
128'h008e00ff00ff00ff020101f3009100ff, /* 2741 */
128'h02008900ff00ff00ff03020201f40201, /* 2742 */
128'h02008500ff00ff00ff03020201f80201, /* 2743 */
128'h018401ff008200ff00ff00ff01fe0201, /* 2744 */
128'hff0201018401ff02010200fd00ff00ff, /* 2745 */
128'h0200f700ff00ff018a01ff00fb00ff00, /* 2746 */
128'h028201e600f400ff00ff018b01ff0201, /* 2747 */
128'h028201e500f100ff00ff019c0282018a, /* 2748 */
128'hff00ff030202019b02010182008a0182, /* 2749 */
128'h020102009203020201e302010200ed00, /* 2750 */
128'h019c009801e4020100eb00ff00ff019b, /* 2751 */
128'h020102009a03020201e400e700ff00ff, /* 2752 */
128'h0201009e020101e400e500ff00ff019a, /* 2753 */
128'h9c00a001e402010200e100ff00ff019b, /* 2754 */
128'h02019a00a201e4020100e000ff00ff01, /* 2755 */
128'h9b00a403020201e400dd00ff00ff0302, /* 2756 */
128'hff019c00a601e600db00ff00ff020101, /* 2757 */
128'h00ff019c02010200a701e600d900ff00, /* 2758 */
128'h00ff019c020100aa020101e600d500ff, /* 2759 */
128'h00ff019d020100aa01e6020100d400ff, /* 2760 */
128'hff00ff019e00ac01e602010200d100ff, /* 2761 */
128'hcd00ff00ff019f00ae020101e700cf00, /* 2762 */
128'h0200cb00ff00ff019f00ae01e7020100, /* 2763 */
128'h01ea00c900ff00ff01a000ae01e80201, /* 2764 */
128'he9020100c700ff00ff030202019f00b0, /* 2765 */
128'h02010200c500ff00ff020101a000b001, /* 2766 */
128'h01eb00c300ff00ff01a1020100b001ea, /* 2767 */
128'h0200c000ff00ff01a202010200b10201, /* 2768 */
128'hbf00ff00ff01a202010200b101eb0201, /* 2769 */
128'hed020100be00ff00ff01a400b201ee00, /* 2770 */
128'h010200bb00ff00ff03020201a300b201, /* 2771 */
128'hb301ef00ba00ff00ff01a600b301ed02, /* 2772 */
128'h0201a600b301f000b800ff00ff01a700, /* 2773 */
128'h00ff01a800b301f100b600ff00ff0302, /* 2774 */
128'h00ff00ff020101a800b201f300b500ff, /* 2775 */
128'h00b200ff00ff01aa00b201f2020100b4, /* 2776 */
128'hff00ff03020201a8020100b201f30201, /* 2777 */
128'h00ff01ab02010200b1020101f400b000, /* 2778 */
128'h00ff00ff020101ac00b001f700ae00ff, /* 2779 */
128'h00ac00ff00ff01ae00b0020101f700ad, /* 2780 */
128'hf900aa00ff00ff03020201ad00b001f8, /* 2781 */
128'hae01fb00a900ff00ff020101af00af01, /* 2782 */
128'hae020101f9020100a800ff00ff01b100, /* 2783 */
128'hb200ac01fd00a700ff00ff020101b000, /* 2784 */
128'h0182020101c500a400ff00ff03020201, /* 2785 */
128'hb4020100aa03020201a602010183008b, /* 2786 */
128'h010182009001c5020100a400ff00ff01, /* 2787 */
128'h0100a200ff00ff01b600aa020101a502, /* 2788 */
128'h0200a701a5020102009603020201c102, /* 2789 */
128'h01a6009a01c300a000ff00ff01b70201, /* 2790 */
128'h009c01c200a000ff00ff020101b800a6, /* 2791 */
128'hc1009e00ff00ff01bb00a403020201a4, /* 2792 */
128'h00ff020101bb00a201a302010200a001, /* 2793 */
128'h0102009f020101a300a301c1009d00ff, /* 2794 */
128'ha500a4020101bf009c00ff00ff01bd02, /* 2795 */
128'h009b00ff00ff03020201bd0201009e01, /* 2796 */
128'h009a00ff00ff01c2009a01a600a601bf, /* 2797 */
128'hff01c3009801a502010200a7020101be, /* 2798 */
128'h01a4020100a901be020102009900ff00, /* 2799 */
128'h9800ff00ff01c4028201010093030202, /* 2800 */
128'h0101ca008b0182020101a800aa01bf00, /* 2801 */
128'h01ac00ab03020201bd009800ff00ff02, /* 2802 */
128'h01ac00ad01be009600ff00ff01cd0088, /* 2803 */
128'hbe009400ff00ff03020201cb02010088, /* 2804 */
128'hff00ff01cd0201008801ab00ae020101, /* 2805 */
128'h0201008801ab00ae03020201bd009400, /* 2806 */
128'h0100b001bd020102009300ff00ff01cd, /* 2807 */
128'h01009200ff00ff01ce0201008801a902, /* 2808 */
128'hff01ce0201008801a9020100b001be02, /* 2809 */
128'hcf0201008801aa00b101be009200ff00, /* 2810 */
128'h01008801aa00b101bf009000ff00ff01, /* 2811 */
128'h02a3019d008e00ff00ff03020201ce02, /* 2812 */
128'hff00ff03020201ce0201008801a900b2, /* 2813 */
128'h8801a8020100d7018202010198008e00, /* 2814 */
128'hda0198008e00ff00ff020101cf020100, /* 2815 */
128'h8c00ff00ff01d10201008801a8020100, /* 2816 */
128'hd10201008801a8020100dc0201019600, /* 2817 */
128'h8801a900dd02010195008c00ff00ff01, /* 2818 */
128'ha900de0195008b00ff00ff01d2020100, /* 2819 */
128'h010194008a00ff00ff01d20201008801, /* 2820 */
128'h8a00ff00ff01d20201008801a900df02, /* 2821 */
128'h01008801a8020100e002010192020100, /* 2822 */
128'ha8020100e10194008800ff00ff01d302, /* 2823 */
128'h910201008800ff00ff01d30201008801, /* 2824 */
128'hff020101d20201008801a900e2020101, /* 2825 */
128'ha202820101008c02010191008800ff00, /* 2826 */
128'h8800ff00ff01d30201008801aa00b101, /* 2827 */
128'haa00b101a4020102008b030202019000, /* 2828 */
128'h010190008600ff00ff01d40201008801, /* 2829 */
128'hd30201008801aa00b101a60201008c02, /* 2830 */
128'ha80201008c0190008600ff00ff020101, /* 2831 */
128'hff00ff01d50201008801a9020100b001, /* 2832 */
128'haa00b001aa008c0201018d0201008500, /* 2833 */
128'h8e008400ff00ff020101d40201008801, /* 2834 */
128'h01008801ab00ae01ab0201008c020101, /* 2835 */
128'hac0201008c018e008400ff00ff01d502, /* 2836 */
128'h8400ff00ff01d50201008801ac00ad01, /* 2837 */
128'h8801ab020100ac01af008c0201018c00, /* 2838 */
128'h018a020102008200ff00ff01d6020100, /* 2839 */
128'h8801ad00aa03020201ae0201008c0201, /* 2840 */
128'h8b0201008300ff00ff020101d4020100, /* 2841 */
128'h01008801ac020100aa01b10201008c01, /* 2842 */
128'h8c020101890201008400ff00ff01d402, /* 2843 */
128'hff020101d20201008801ae00a801b400, /* 2844 */
128'ha701b40201008c02010189008500ff00, /* 2845 */
128'h8500ff00ff020101d10201008801af00, /* 2846 */
128'h01b000a403020201b50201008c018a00, /* 2847 */
128'h02010188008600ff00ff01d102010088, /* 2848 */
128'h0201008801af020100a4020101b8008c, /* 2849 */
128'h0201008c0188008700ff00ff020101cf, /* 2850 */
128'h00ff00ff01cf0201008801b200a101ba, /* 2851 */
128'h008801b3009e01be008c020101860088, /* 2852 */
128'h02010185008900ff00ff020101cd0201, /* 2853 */
128'h0201008801b30201009c01bf0201008c, /* 2854 */
128'h0201008c0185008a00ff00ff020101cc, /* 2855 */
128'h00ff00ff01cc0201008801b7009701c2, /* 2856 */
128'h008801b8009401c6008c02010184008a, /* 2857 */
128'h018300fd00ff0101008c020101ca0201, /* 2858 */
128'h0101008e0182020101c60201008c0201, /* 2859 */
128'h0202008c020101c90201008801b80282, /* 2860 */
128'h8a028201ca0201008c018300fd00ff03, /* 2861 */
128'h830201008c01c90201008801bb028201, /* 2862 */
128'h01bf028601d0008c02010200fc00ff01, /* 2863 */
128'h00fb00ff0185008c020101c702010088, /* 2864 */
128'hc602010088019601ff0201008c020102, /* 2865 */
128'h8c010100fb00ff01850201008c020101, /* 2866 */
128'h01008c01c602010088019701ff020100, /* 2867 */
128'h010088019901ff008800ff00ff018602, /* 2868 */
128'h01008700ff00ff0188008c020101c402, /* 2869 */
128'h880201008c01c402010088019901ff02, /* 2870 */
128'hc202010088019b01ff008600ff00ff01, /* 2871 */
128'hff0201008500ff00ff018a008c020101, /* 2872 */
128'h8a0201008c020101c102010088019b01, /* 2873 */
128'h010089019b01ff0201008400ff00ff01, /* 2874 */
128'hff008300ff00ff018b0201008c01c102, /* 2875 */
128'hff00ff018d008c020101c00089019d01, /* 2876 */
128'h0101bf008a0201019b01ff0201008200, /* 2877 */
128'h8601b2020100ff00ff018e0201008c02, /* 2878 */
128'hff018f0201008c01c0008a020101e202, /* 2879 */
128'hbe008a01e002820188028201b100fe00, /* 2880 */
128'h8f01b0020100fd00ff0191008c020101, /* 2881 */
128'h01910201008c01bd020102008b01dc00, /* 2882 */
128'h0101d5020102009601ad020100fc00ff, /* 2883 */
128'hfb00ff01920201008c01bd0201008c02, /* 2884 */
128'h03020201d3020102009803020201ac00, /* 2885 */
128'h020100fa00ff0194008c020101bd008b, /* 2886 */
128'h0201008c020101bd008c01d3009c01ac, /* 2887 */
128'hcf0201009f03020201ab00f900ff0194, /* 2888 */
128'h95020102008b03020201bb0201008c01, /* 2889 */
128'h020201cc02010200a001ac00f900ff01, /* 2890 */
128'hf900ff01960201008c020101bd008b03, /* 2891 */
128'h8c01be008c020101ca020100a401aa00, /* 2892 */
128'h8b01cc00a401aa00f800ff0198020100, /* 2893 */
128'h00f800ff019a008c020101bb02010200, /* 2894 */
128'h01008c01be008b01c802010200a601a9, /* 2895 */
128'h8c020101c500a901a800f800ff019a02, /* 2896 */
128'ha700f800ff019b0201008c01bd020100, /* 2897 */
128'h008c020101bd008b03020201c400aa01, /* 2898 */
128'h01bd008c01c300ab01a700f800ff019d, /* 2899 */
128'h00ac01a600f800ff019d0201008c0201, /* 2900 */
128'h01008c03020201bb0201008c020101c1, /* 2901 */
128'h01be02010200ad01a500f800ff019e02, /* 2902 */
128'hf800ff01a0008c020101bd008b030202, /* 2903 */
128'h0101bd008c020101be00ae020101a400, /* 2904 */
128'h03020201a300f900ff019f0201008c02, /* 2905 */
128'h008c01bd0201008c020101bb020100af, /* 2906 */
128'h01bc020100b001a400f900ff01a00201, /* 2907 */
128'h00b001a400f900ff01a2008c01be008b, /* 2908 */
128'h01a20201008c020101bd008c020101ba, /* 2909 */
128'hbb020102008b01bb00b101a300f900ff, /* 2910 */
128'h020101a200f900ff01a4008b03020201, /* 2911 */
128'h01a40201008c020101bd008b01b900b2, /* 2912 */
128'h01be008c020101b600b201a200fa00ff, /* 2913 */
128'h01b500b201a200fa00ff01a50201008c, /* 2914 */
128'h01a7008c020101bb020102008b030202, /* 2915 */
128'h008c020101b400b201a1020100fa00ff, /* 2916 */
128'h020100fa00ff01a70201008c020101bd, /* 2917 */
128'h0201008c01bd0201008c01b400b201a1, /* 2918 */
128'h008b01b400b201a1020100fb00ff01a7, /* 2919 */
128'h00b201a1020100fb00ff01a9008c01be, /* 2920 */
128'h01a90201008c020101bd008c020101b1, /* 2921 */
128'h0201008c020101b000b201a200fb00ff, /* 2922 */
128'h00b201a200fb00ff01aa0201008c01bd, /* 2923 */
128'h00fb00ff01ac008c020101bd008b01b1, /* 2924 */
128'h03020201bc008c01af00b201a0020102, /* 2925 */
128'h9f02010200fb00ff020101ab0201008c, /* 2926 */
128'h020201bb020102008b01af00b2020101, /* 2927 */
128'h0201ac00b201a200fb00ff01ae008b03, /* 2928 */
128'h00fc00ff01af008c020101bd008b0302, /* 2929 */
128'h01ae0201008c01be008c01ad00b001a2, /* 2930 */
128'hbc020102008b01ad00b001a200fd00ff, /* 2931 */
128'h00af03020201a100fd00ff01b0008c01, /* 2932 */
128'h01af0201008c020101bd008b01ab0201, /* 2933 */
128'h008c01ab00ae020101a100fe00ff0201, /* 2934 */
128'h00fe00ff020101b00201008c01bd0201, /* 2935 */
128'h008c020101bd008b01ab00ae020101a1, /* 2936 */
128'h020101a900ac01a300fe00ff020101b2, /* 2937 */
128'hfe00ff03020201b10201008c01be008c, /* 2938 */
128'hbd0201008c020101a800ab01a3020100, /* 2939 */
128'h01a400fe00ff03020201b20201008c01, /* 2940 */
128'hb5008c020101bd008b03020201a800aa, /* 2941 */
128'h0101bd008c01a800aa01a400ff00ff01, /* 2942 */
128'ha901a2000100ff00ff01b50201008c02, /* 2943 */
128'h01b50201008c01be008c01a702010200, /* 2944 */
128'h020100aa0201019f0201008200ff00ff, /* 2945 */
128'hff01b7008c020101bd008b03020201a6, /* 2946 */
128'hbd008c01a800aa019f0201008200ff00, /* 2947 */
128'h8200ff00ff020101b60201008c020101, /* 2948 */
128'h0102008b01a900aa0201019c02010200, /* 2949 */
128'h008200ff00ff01b9008b03020201bb02, /* 2950 */
128'h03020201a6020100aa0201019b020102, /* 2951 */
128'h00ff00ff01b90201008c028201bc008b, /* 2952 */
128'h008c020101a8009c0101008c019c0083, /* 2953 */
128'h019a008400ff00ff01b90201008c01be, /* 2954 */
128'h008b03020201a8009a030202008d0201, /* 2955 */
128'h8500ff00ff01bb008c020101bb020102, /* 2956 */
128'ha802010200960184020102008c019900, /* 2957 */
128'hff020101ba0201008c020101bd008c01, /* 2958 */
128'h020102008f018b008c0198008500ff00, /* 2959 */
128'hff03020201ba0201008c01be008c01aa, /* 2960 */
128'h820201018a008d02010196008500ff00, /* 2961 */
128'h01bd008b03020201aa02010182008a01, /* 2962 */
128'h0195008600ff00ff020101bc008c0201, /* 2963 */
128'hbd008c01ae0287018f020102008c0201, /* 2964 */
128'h94008700ff00ff01bd0201008c020101, /* 2965 */
128'hff01bd0201008c01be008c01c6008c01, /* 2966 */
128'h0201c4008d020101910201008800ff00, /* 2967 */
128'h00ff020101be008c020101bd008b0302, /* 2968 */
128'h0101c5008c0201018f020102008800ff, /* 2969 */
128'hff00ff01bf0201008c020101bd008c02, /* 2970 */
128'h01c50201008c030202018e0201008900, /* 2971 */
128'h00ff01c1008b03020201bb020102008b, /* 2972 */
128'h020101bd008b01c7008c018f008900ff, /* 2973 */
128'h008c018c0201008b00ff00ff01c1008c, /* 2974 */
128'h00ff01c10201008c01be008c020101c5, /* 2975 */
128'h008b01c6008d0201018a0201008b00ff, /* 2976 */
128'h8b00ff00ff01c3008c020101bb020102, /* 2977 */
128'h01bd008b01c5020102008c0201018a00, /* 2978 */
128'h0189008d00ff00ff01c20201008c0201, /* 2979 */
128'h00ff01c20201008c01be008c01c6008c, /* 2980 */
128'h8b03020201c4008d02010187008e00ff, /* 2981 */
128'h8e00ff00ff020101c3008c020101bd00, /* 2982 */
128'h0101bd008c020101c5008c0201018600, /* 2983 */
128'h8c0185008f00ff00ff01c40201008c02, /* 2984 */
128'hff01c40201008c01bd0201008c01c600, /* 2985 */
128'h008b03020201c4008d0183009100ff00, /* 2986 */
128'h0282009100ff00ff01c6008c020101bd, /* 2987 */
128'h0201008c020101bd008c020101c5008c, /* 2988 */
128'h008b01c6008c0182009200ff00ff01c5, /* 2989 */
128'h00ff00ff01c7008b03020201bb020102, /* 2990 */
128'h01c7008c020101bd008b01c50201009f, /* 2991 */
128'h008c020101bd008c01c6009e00ff00ff, /* 2992 */
128'h008b01c6009e00ff00ff020101c60201, /* 2993 */
128'hc5009c00ff00ff01c9008b03020201bd, /* 2994 */
128'h01c80201008c020101bd008b03020201, /* 2995 */
128'h0101028301a7008c01c6009c00ff00ff, /* 2996 */
128'h00ff00ff020101c70201008c01900283, /* 2997 */
128'h01018e008701a6020102008b01c6009d, /* 2998 */
128'h03020201c5009b00ff00ff01ca008c02, /* 2999 */
128'h01018602010200910182020101a1008b, /* 3000 */
128'h0101c5009b00ff00ff01c90201008c02, /* 3001 */
128'h018402010097030202019f0201008c02, /* 3002 */
128'h008b01c6009b00ff00ff01ca0201008c, /* 3003 */
128'hff01cc008c04030203009903020201a0, /* 3004 */
128'hcb020100a901a1008c01c3009c00ff00, /* 3005 */
128'h9e0201008c020101c1009d00ff00ff01, /* 3006 */
128'h9f00ff00ff020101ca020100aa020101, /* 3007 */
128'ha9030202019f008b03020201be020100, /* 3008 */
128'haa01a0008c01be00a000ff00ff01cd00, /* 3009 */
128'h8b01bd020100a100ff00ff01cc020100, /* 3010 */
128'hff00ff01ce00a9030202019d02010200, /* 3011 */
128'hff01ce00aa0201019f008b01bc00a200, /* 3012 */
128'h0100a901a1008c020101b900a300ff00, /* 3013 */
128'h02008b01b900a500ff00ff020101cc02, /* 3014 */
128'hff00ff03020201cc00aa0201019e0201, /* 3015 */
128'h00ab03020201a0008b01b6020100a600, /* 3016 */
128'h8c020101b202010200a800ff00ff01cb, /* 3017 */
128'hb200a900ff00ff01c9020100ad01a200, /* 3018 */
128'hff01c900ae01a0020102008b03020201, /* 3019 */
128'hff01c900ae01a3008c01b100ab00ff00, /* 3020 */
128'hc600b001a20201008c01af00ac00ff00, /* 3021 */
128'h01a4008b03020201ad00ae00ff00ff01, /* 3022 */
128'h020101ab00af00ff00ff020101c500b0, /* 3023 */
128'h00ff00ff020101c400b0020101a4008c, /* 3024 */
128'hc500b001a4020102008b01aa020100b1, /* 3025 */
128'h03020201a5008b01a900b200ff00ff01, /* 3026 */
128'h0101a402010200b300ff00ff01c300b1, /* 3027 */
128'hb500ff00ff01c200b2020101a6008c02, /* 3028 */
128'h00ff01c200b201a6020102008b01a600, /* 3029 */
128'h020201be00b301a9008b01a400b600ff, /* 3030 */
128'hb301aa008c01a0020100b800ff00ff03, /* 3031 */
128'h008b019f02010200ba00ff00ff01be00, /* 3032 */
128'h9c00bc00ff00ff01be00b301a9020102, /* 3033 */
128'h00ff020101bc00b301ac008b03020201, /* 3034 */
128'h01bc00b301ac0201008c019b00be00ff, /* 3035 */
128'h01bb00b201ae008b019b00bf00ff00ff, /* 3036 */
128'h008c02010195020100c200ff00ff0201, /* 3037 */
128'h9400c400ff00ff01bb00b103020201ae, /* 3038 */
128'h01ba00b103020201ae0201008c020101, /* 3039 */
128'h01b900b001b2008b019400c600ff00ff, /* 3040 */
128'h01b2008c0201019100c700ff00ff0201, /* 3041 */
128'h8f02010200c900ff00ff01b900b00201, /* 3042 */
128'h00ff020101b700b001b2020102008b01, /* 3043 */
128'hb600af01b6008b030202018c00cc00ff, /* 3044 */
128'hae01b7008c018b00ce00ff00ff020101, /* 3045 */
128'h008b018902010200cf00ff00ff01b700, /* 3046 */
128'h0100d200ff00ff01b600ae01b6020102, /* 3047 */
128'h020201b300ad01ba008b030202018502, /* 3048 */
128'hba008c02010183020100d400ff00ff03, /* 3049 */
128'hff00ff020101b202010200aa03020201, /* 3050 */
128'h00aa020101ba020102008b018400d700, /* 3051 */
128'h00a801bf008c010100d800ff00ff01b5, /* 3052 */
128'h01b200a601c0020100e500ff00ff01b5, /* 3053 */
128'h00a503020201c100e600ff00ff030202, /* 3054 */
128'h020100a301c500e600ff00ff01b20201, /* 3055 */
128'h03020201c302010200e700ff00ff01b1, /* 3056 */
128'h01b3009e01c900e600ff00ff01b300a1, /* 3057 */
128'hff01b3009a03020201c900e800ff00ff, /* 3058 */
128'haf020102009903020201c900eb00ff00, /* 3059 */
128'h0201b2009401cb00ee00ff00ff020101, /* 3060 */
128'h008d0101028201cb00f000ff00ff0302, /* 3061 */
128'h020100f400ff00ff03020201b1020102, /* 3062 */
128'h020201b20201018400840184020101ca, /* 3063 */
128'hfb00ff00ff018a01ff00f700ff00ff03, /* 3064 */
128'hfe00ff00ff030202018201ff02010200, /* 3065 */
128'h8200ff00ff00ff03020201ff02010200, /* 3066 */
128'h01fd008500ff00ff00ff03020201fd00, /* 3067 */
128'hff00ff03020201f5008900ff00ff00ff, /* 3068 */
128'hff00ff00ff01f102010182008d00ff00, /* 3069 */
128'h009600ff00ff00ff01ee020102009100, /* 3070 */
128'h020102009c00ff00ff00ff01e8020102, /* 3071 */
128'h0201de020102009f00ff00ff00ff01e3, /* 3072 */
128'h01d70282010100a400ff00ff00ff0302, /* 3073 */
128'hff00ff01d500ab00ff00ff00ff030202, /* 3074 */
128'hff0182020101cb0201018200b000ff00, /* 3075 */
128'h82028201c20201018300b500ff00ff00, /* 3076 */
128'h0201bb0201018200be00ff00ff00ff01, /* 3077 */
128'h00ff00ff01bb00c600ff00ff00ff0302, /* 3078 */
128'h00ff0184028301a20283018400cd00ff, /* 3079 */
128'h0185028401980284018400d700ff00ff, /* 3080 */
128'h00ff00ff00ff019100e600ff00ff00ff, /* 3081 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3082 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3083 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3084 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3085 */
128'h00a800ff00ff00ff00ff00ff00ff00ff, /* 3086 */
128'h00ff00ff059500f100ff00ff00ff058e, /* 3087 */
128'h059600ed00ff00ff00ff059500ee00ff, /* 3088 */
128'h00ff00ff00ff059600ed00ff00ff00ff, /* 3089 */
128'h00ff059600ed00ff00ff00ff059600ed, /* 3090 */
128'h00ff0596009e058600d8058500eb00ff, /* 3091 */
128'h05960094059900c4059900f3058e00e0, /* 3092 */
128'h00bd05a000a4059600b005a200d200ff, /* 3093 */
128'h059800a805b200c800ff05960091059f, /* 3094 */
128'h00c800ff0596008d05a700b505a700a1, /* 3095 */
128'h008b05ab00b105aa00a0059800a505b5, /* 3096 */
128'h05b0009d059900a105b800c800ff0596, /* 3097 */
128'h009f05ba00c800ff0596008805b000ac, /* 3098 */
128'h00ff0596008605b600a505b5009b0599, /* 3099 */
128'h05b700a505b6009a0599009d05bc00c8, /* 3100 */
128'h00990599009b05be00c800ff05960085, /* 3101 */
128'h05bf00c800ff0596008305bc00a005b9, /* 3102 */
128'h0596008205be009e05bb00980599009a, /* 3103 */
128'h009d05bd00960599009905c000c800ff, /* 3104 */
128'h0599009705c200c800ff0596008205bf, /* 3105 */
128'h00c800ff0596008205c1009c05bc0096, /* 3106 */
128'h008205c2009b05bd00950599009605c3, /* 3107 */
128'h05be00940599009505c400c800ff0596, /* 3108 */
128'h009505c400c800ff0596008305c2009a, /* 3109 */
128'h00ff0596008305c3009905bf00930599, /* 3110 */
128'h05c4009905bf0091059a009405c500c8, /* 3111 */
128'h0091059a009405c500c800ff05960083, /* 3112 */
128'h05c700c800ff0596008305c5009805bf, /* 3113 */
128'h0596008405c5009805be0091059a0092, /* 3114 */
128'h009805bf0090059a009205c700c800ff, /* 3115 */
128'h059a009205c700c800ff0596008505c4, /* 3116 */
128'h00c800ff0596008505c5009705c0008f, /* 3117 */
128'h008505c6009705bf008f059a009105c8, /* 3118 */
128'h05be008f059a009105c800c800ff0596, /* 3119 */
128'h009105c800c800ff0596008605c50098, /* 3120 */
128'h008605c600970592008f059d008f059a, /* 3121 */
128'h059a009005a00090059900c800ff0596, /* 3122 */
128'h0596008905a80097058d0096059b008e, /* 3123 */
128'h0090059e0092059900c800ff05960086, /* 3124 */
128'h008e05a60097058b0099059a008e059a, /* 3125 */
128'h059c0094059900c800ff059600870592, /* 3126 */
128'h05a300960587009e0599008e059a0090, /* 3127 */
128'h0096059a00c700ff05960088058d0096, /* 3128 */
128'h0098058200a20599008d059a008f059b, /* 3129 */
128'h059a00c700ff059600880589009c05a1, /* 3130 */
128'h050100a30599008d059a008f059b0096, /* 3131 */
128'h00c700ff059600890587009e05a10097, /* 3132 */
128'h00ba0599008d059a008f059a0097059a, /* 3133 */
128'h009f058400e40596008a058300a305a0, /* 3134 */
128'h008f05990098059a00990585009a0587, /* 3135 */
128'h008a058300a4059f00ba0599008d059a, /* 3136 */
128'h009905910096058b00aa058e00a50596, /* 3137 */
128'h008d059a008f05990098059a0093058b, /* 3138 */
128'h009f059800a1059500b2059e00ba0599, /* 3139 */
128'h0098059a008e05900099059300940591, /* 3140 */
128'h00b3059e00b90599008d059a008f0599, /* 3141 */
128'h0098059400930595009a059b00a00595, /* 3142 */
128'h008d059a008f05990098059a008c0592, /* 3143 */
128'h009705a1009d059500b4059d00b90599, /* 3144 */
128'h0098059a008905960097059400930595, /* 3145 */
128'h00b5059c00b7059b008d059a008f0599, /* 3146 */
128'h0096059400930596009505a5009b0595, /* 3147 */
128'h008e059a008f05980099059a00890596, /* 3148 */
128'h009405a7009a059500b5059c00b6059b, /* 3149 */
128'h0099059a008905960096059400930596, /* 3150 */
128'h00b6059b00b5059c008e059a008f0598, /* 3151 */
128'h0095059400930596009305aa00980595, /* 3152 */
128'h008e059a008f05980099059a008a0596, /* 3153 */
128'h009305ac0096059500b7059b00b1059f, /* 3154 */
128'h0098059a008a05960095059300940596, /* 3155 */
128'h00b7059b00ad05a3008e059a008f0599, /* 3156 */
128'h0094059400940596009305ac00960595, /* 3157 */
128'h008f059a008f05990098059a008b0595, /* 3158 */
128'h009505ac0095059500b7059c00a905a5, /* 3159 */
128'h0098059a008b05960093059400930596, /* 3160 */
128'h00b8059b00a405aa008f059a008f0599, /* 3161 */
128'h0093059400930596009705ac00930595, /* 3162 */
128'h008f059a008f05990098059a008b0596, /* 3163 */
128'h009705ac0093059500b8059b00a005ae, /* 3164 */
128'h0097059a008b05960093059300940596, /* 3165 */
128'h00b8059b009e05b0008f059a008f059a, /* 3166 */
128'h0091059500930596009805ac00920595, /* 3167 */
128'h0090059a008f059b0096059a008c0596, /* 3168 */
128'h008b05ac0091059500b9059a009b05b2, /* 3169 */
128'h008c05960091059500920597008d0501, /* 3170 */
128'h009905b40090059a0090059a0096059a, /* 3171 */
128'h008d0583008b05ac0090059500b9059a, /* 3172 */
128'h0095059a008d05950090059600920596, /* 3173 */
128'h00b9059a009705b50091059a0090059b, /* 3174 */
128'h00900597008c0586008b05aa00900595, /* 3175 */
128'h0091059d0092059a008d059500900597, /* 3176 */
128'h008f059500ba0599009505b70091059a, /* 3177 */
128'h0090059700900596008d0586008b05ab, /* 3178 */
128'h0092059a0091059f0090059a008d0595, /* 3179 */
128'h008b05aa008f059500ba0599009405b7, /* 3180 */
128'h008e0595008f059700900596008c0588, /* 3181 */
128'h00ba0599009205b90092059a009105c9, /* 3182 */
128'h00900596008c058a008b05a9008e0595, /* 3183 */
128'h0094059a009205c8008e0596008e0597, /* 3184 */
128'h0088059b008e059500ba0599009105b8, /* 3185 */
128'h008d0599008f0596008b058b008b0586, /* 3186 */
128'h009005b90094059a009205c8008e0596, /* 3187 */
128'h008b0582008e0599008d059500ba0599, /* 3188 */
128'h008e0596008d059a008e0595008c058c, /* 3189 */
128'h00ba0599008f05b90095059a009205c8, /* 3190 */
128'h008d0596008b058f009b0597008d0595, /* 3191 */
128'h0097059a009305c7008f0595008d059a, /* 3192 */
128'h009c0597008c059500ba0599008e05b8, /* 3193 */
128'h008f0595008d059a008d0595008c058f, /* 3194 */
128'h00ba0599008d05b90097059a009405c6, /* 3195 */
128'h008c0595008c0590009d0595008c0595, /* 3196 */
128'h0099059a009505c500900595008b059c, /* 3197 */
128'h009c0595008c059500ba0599008c05b8, /* 3198 */
128'h00900595008b059c008c0595008b0592, /* 3199 */
128'h00ba0599008c05b7009a059a009505c5, /* 3200 */
128'h008b0595008b0593009c0594008c0595, /* 3201 */
128'h009d059a009605c400900596008a059d, /* 3202 */
128'h009c0594008b059500ba0599008b05b5, /* 3203 */
128'h009105950089059e008a0596008b0594, /* 3204 */
128'h00b9059a008b05b3009f059a009705c3, /* 3205 */
128'h008a0595008c0593009d0594008b0595, /* 3206 */
128'h00a0059a009905c1009105950089059e, /* 3207 */
128'h009e0593008b059500b9059a008a05b3, /* 3208 */
128'h009105950089059f00880596008c0593, /* 3209 */
128'h00b9059a008a05ae00a5059a009a05c0, /* 3210 */
128'h00880596008b0593009f0593008b0595, /* 3211 */
128'h00aa059a009c05be009105960088059f, /* 3212 */
128'h00a00592008b059500b8059b008905aa, /* 3213 */
128'h00920595008705a000880596008b0593, /* 3214 */
128'h00b8059b008905a800ac059a009d05bd, /* 3215 */
128'h00870595008c059200a10593008a0595, /* 3216 */
128'h00b1059a009f05bb00920595008705a1, /* 3217 */
128'h00a10593008a059500b8059b008905a3, /* 3218 */
128'h00930594008605a200870595008c0592, /* 3219 */
128'h00b8059a008a05a000b4059a009f05bb, /* 3220 */
128'h00860594008d059200a10593008a0595, /* 3221 */
128'h00b6059a009f05bb00930595008505a3, /* 3222 */
128'h00a10593008b059400b7059b008a059e, /* 3223 */
128'h00930595008505a300850595008d0592, /* 3224 */
128'h00b7059b0089059d00b8059a009e05bc, /* 3225 */
128'h00850595008d059200a10593008b0594, /* 3226 */
128'h00b9059a009d05bd00930596008405a3, /* 3227 */
128'h00a10593008b059400b7059b0089059c, /* 3228 */
128'h00940595008405a400840595008d0592, /* 3229 */
128'h008a059c00b9059a009d059b00890599, /* 3230 */
128'h008d059200a10592008c059400b6059b, /* 3231 */
128'h00940595008305920001059200830596, /* 3232 */
128'h008a059a00bb059a009c059c00890599, /* 3233 */
128'h008e059200a10592008c059400b5059c, /* 3234 */
128'h00940595008305920001059200830595, /* 3235 */
128'h008a059a00bb059a009b059c008a0599, /* 3236 */
128'h008e059300a00592008c059400b5059c, /* 3237 */
128'h00950595008205920082059200820595, /* 3238 */
128'h00a605010094059a009a059c008b0599, /* 3239 */
128'h009f0593008c059400b4059d008a059a, /* 3240 */
128'h008205910083059200820595008e0593, /* 3241 */
128'h0093059a0099059c008c059900950595, /* 3242 */
128'h008b058300a5059d008b059a00a40584, /* 3243 */
128'h00820595008f0592009f0593008c0594, /* 3244 */
128'h008c0599009605940082059100830592, /* 3245 */
128'h008b059a00a305850093059a0099059c, /* 3246 */
128'h009e0592008d0594008b058400a3059e, /* 3247 */
128'h0096059400010592008305a800900593, /* 3248 */
128'h00a105880092059a0098059c008d0599, /* 3249 */
128'h008d0594008a058700a0059f008b059a, /* 3250 */
128'h009605a7008405a700900593009d0593, /* 3251 */
128'h009e058a0092059a0097059c008e0599, /* 3252 */
128'h008d05940089058a009c05a0008d059a, /* 3253 */
128'h009605a6008605a500910594009c0593, /* 3254 */
128'h009c058c0091059a0097059c008e0599, /* 3255 */
128'h008d05940088058d009905a1008d059b, /* 3256 */
128'h009705a5008605a500910595009a0594, /* 3257 */
128'h0099058f0091059a0095059d008f0599, /* 3258 */
128'h008d05940088058f009505a2008e059b, /* 3259 */
128'h009805a3008705a50092059500980595, /* 3260 */
128'h009405920091059a0095059c00900599, /* 3261 */
128'h008e059400870594008e05a5008e059d, /* 3262 */
128'h009805a3008705a50092059500970595, /* 3263 */
128'h009005950090059a0094059c00910599, /* 3264 */
128'h008e059400860599008605a8008f059f, /* 3265 */
128'h009805a3008805a30094059600940596, /* 3266 */
128'h009005c4009005990094059c00910599, /* 3267 */
128'h0094059700910598008e0594008605c7, /* 3268 */
128'h0093059c00920599009805a3008805a3, /* 3269 */
128'h008f0594008505c8009005c400900599, /* 3270 */
128'h009905a2008805a300940599008e0598, /* 3271 */
128'h009205c3009005990092059c00930599, /* 3272 */
128'h0095059d0084059c00900594008505c7, /* 3273 */
128'h0091059c00940599009905a1008a05a2, /* 3274 */
128'h00900594008405c7009305c300900599, /* 3275 */
128'h00950598009905a1008a05a2009505bd, /* 3276 */
128'h008305c8009405c3008f05990091059c, /* 3277 */
128'h009a05a0008b05a0009705bc00900594, /* 3278 */
128'h009505c3008f05990091059b00950599, /* 3279 */
128'h008b05a0009805ba00910594008305c7, /* 3280 */
128'h008e0599008f059c00970598009a05a0, /* 3281 */
128'h009905ba00910594008205c7009705c3, /* 3282 */
128'h008f059c00970598009b059e008c059f, /* 3283 */
128'h00930594008205c6009905c2008e0599, /* 3284 */
128'h00980598009b059e008d059e009a05b7, /* 3285 */
128'h008205c5009b05c1008e0599008e059c, /* 3286 */
128'h009b059d008e059e009b05b600930594, /* 3287 */
128'h009d05c0008e0599008e059b00990598, /* 3288 */
128'h008e059e009c05b400940594008205c4, /* 3289 */
128'h008e0599008d059c00990598009c059c, /* 3290 */
128'h009e05b200950594008205c4009d05c0, /* 3291 */
128'h008c059c009a0598009c059c008f059c, /* 3292 */
128'h00960594008305c200a005bd008f0599, /* 3293 */
128'h009a0598009c059c008f059c009f05b0, /* 3294 */
128'h008405bf00a305bb00900599008c059c, /* 3295 */
128'h009c059b0091059a00a105ae00970594, /* 3296 */
128'h00a505b800920599008c059b009b0598, /* 3297 */
128'h0091059a00a305aa00990594008605bc, /* 3298 */
128'h00950599008c059a009c0598009d059a, /* 3299 */
128'h00a305aa00990594008705b900a905b3, /* 3300 */
128'h008e0597009d0598009e059900920599, /* 3301 */
128'h009b0594008805b800aa05b100960599, /* 3302 */
128'h009d0598009e05990092059900a505a6, /* 3303 */
128'h008b05b300ae05ac0099059900900595, /* 3304 */
128'h009e05980093059800a805a1009e0594, /* 3305 */
128'h00b305a6009c059900920592009e0598, /* 3306 */
128'h0094059700aa059e009f0594008d05af, /* 3307 */
128'h009f05990094058f009f0598009e0598, /* 3308 */
128'h00ad059800a20594008e05ac00b705a1, /* 3309 */
128'h0097058c009f0598009f059600950597, /* 3310 */
128'h00a70591009405a600bf059700a40599, /* 3311 */
128'h009c058800d70592009a059200b6058e, /* 3312 */
128'h00a5058700c3058700d4059e00fe0596, /* 3313 */
128'h0599008800ff058800a6058600da0586, /* 3314 */
128'h00ff00ff00ff058b00f100ff00ff00ff, /* 3315 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3316 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3317 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3318 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3319 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3320 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3321 */
128'h00ff00ff00ff00ff00ff00ff00ff00ff, /* 3322 */
128'h009b058600e300ff00ff00ff00ff00ff, /* 3323 */
128'h00af0585008505840097058b009a0589, /* 3324 */
128'h008605840096058c00b305870099058c, /* 3325 */
128'h009b0586009d058600b5058a00980583, /* 3326 */
128'h0098058b009905890085058b009a0589, /* 3327 */
128'h0098058c00af0585008405850097058b, /* 3328 */
128'h00970583008505850096058c00b20589, /* 3329 */
128'h0099058a009a0589009a058800b3058c, /* 3330 */
128'h0097058b0097058c0098058c0083058b, /* 3331 */
128'h00b0058c0097058c00af058500840585, /* 3332 */
128'h00b1058b00980583008505850096058c, /* 3333 */
128'h0082058b0097058c0098058d0097058b, /* 3334 */
128'h0097058b0096058d0097058600010587, /* 3335 */
128'h000105860096058c00af058500830586, /* 3336 */
128'h00980583008505850096058c00af0587, /* 3337 */
128'h00980586000105870097058b00b0058b, /* 3338 */
128'h00970585008405850082058b0097058c, /* 3339 */
128'h00820587009e05840096058500830585, /* 3340 */
128'h00b3058500840585009a058400b30585, /* 3341 */
128'h00b705840098058300850585009a0584, /* 3342 */
128'h00970585008505850097058200840585, /* 3343 */
128'h00870584008905840097058400840584, /* 3344 */
128'h009e0584009605840084058500960584, /* 3345 */
128'h008705840099058400b3058500010588, /* 3346 */
128'h0098058300850585009a058400b30584, /* 3347 */
128'h0097058400870584009e058400b70584, /* 3348 */
128'h00880584008805840097058300850584, /* 3349 */
128'h0097058b009605840084058500960584, /* 3350 */
128'h00b20584008805840099058400b3058e, /* 3351 */
128'h009f058300b1058a0098058d009a0584, /* 3352 */
128'h00970584008405840096058500870584, /* 3353 */
128'h0083058500960584008805840001058b, /* 3354 */
128'h0099058400b3058e0097058b00960585, /* 3355 */
128'h0098058d009a058400b2058400880584, /* 3356 */
128'h0096058500870584009f058300b1058a, /* 3357 */
128'h00960584008805840001058b0097058c, /* 3358 */
128'h00b30588000105850097058b0097058c, /* 3359 */
128'h009a058400b205840088058400990584, /* 3360 */
128'h00870584009f058300b1058a0098058d, /* 3361 */
128'h008805840001058b0098058b00960585, /* 3362 */
128'h00010585009e05840097058c00960584, /* 3363 */
128'h00b30584008705840099058400b30588, /* 3364 */
128'h009e058400b705840098058d009a0584, /* 3365 */
128'h008805850099058a0096058500870584, /* 3366 */
128'h009e05840099058a0097058400860584, /* 3367 */
128'h00860584009a058400b3058700820585, /* 3368 */
128'h0098058300850585009a058400b30584, /* 3369 */
128'h00850585009705010086058400b70584, /* 3370 */
128'h00890584009905840082058400970585, /* 3371 */
128'h008305850096058c009e05850097058e, /* 3372 */
128'h009a058400b3058e009a058400b30586, /* 3373 */
128'h0097058c00b0058b0098058300850585, /* 3374 */
128'h0083058b00980585008205840098058d, /* 3375 */
128'h008305850096058c009e05850097058d, /* 3376 */
128'h009a058400b4058d009a058400b30586, /* 3377 */
128'h0097058b00b1058b0098058300850585, /* 3378 */
128'h0084058b00970585008305840098058d, /* 3379 */
128'h008405850096058c009e05850099058a, /* 3380 */
128'h009a058400b5058a009c058400b30585, /* 3381 */
128'h0098058a00b2058b0098058300850585, /* 3382 */
128'h0086058b0097058400840584009a058a, /* 3383 */
128'h008705830098058a00a00583009c0586, /* 3384 */
128'h009a058300b80586009e058400b40582, /* 3385 */
128'h009d058600b5058a0098058300860584, /* 3386 */
128'h0001058a0098058300850583009d0585, /* 3387 */
128'h00e0354f00e9374f00e0354f0020272d, /* 3388 */
128'hffffca8cffffca7800e1e6e800e9374f, /* 3389 */
128'hffffca8affffcab4ffffca8affffcaa0, /* 3390 */
128'h000000000000000000000000ffffcac6, /* 3391 */
128'he00600003800000039080000edfe0dd0, /* 3392 */
128'h00000000100000001100000028000000, /* 3393 */
128'h0000000000000000a806000059010000, /* 3394 */
128'h00000000010000000000000000000000, /* 3395 */
128'h02000000000000000400000003000000, /* 3396 */
128'h020000000f0000000400000003000000, /* 3397 */
128'h2c6874651b0000001400000003000000, /* 3398 */
128'h007665642d657261622d656e61697261, /* 3399 */
128'h2c687465260000001000000003000000, /* 3400 */
128'h0100000000657261622d656e61697261, /* 3401 */
128'h1a0000000300000000006e65736f6863, /* 3402 */
128'h313440747261752f636f732f2c000000, /* 3403 */
128'h0000003030323531313a303030303030, /* 3404 */
128'h00000000737570630100000002000000, /* 3405 */
128'h01000000000000000400000003000000, /* 3406 */
128'h000000000f0000000400000003000000, /* 3407 */
128'h20a10700380000000400000003000000, /* 3408 */
128'h03000000000000304075706301000000, /* 3409 */
128'h0300000080f0fa024b00000004000000, /* 3410 */
128'h03000000007570635b00000004000000, /* 3411 */
128'h03000000000000006700000004000000, /* 3412 */
128'h0000000079616b6f6b00000005000000, /* 3413 */
128'h7a6874651b0000001300000003000000, /* 3414 */
128'h0000766373697200656e61697261202c, /* 3415 */
128'h34367672720000000b00000003000000, /* 3416 */
128'h0b000000030000000000636466616d69, /* 3417 */
128'h0000393376732c76637369727c000000, /* 3418 */
128'h01000000850000000000000003000000, /* 3419 */
128'h6f72746e6f632d747075727265746e69, /* 3420 */
128'h04000000030000000000000072656c6c, /* 3421 */
128'h0000000003000000010000008f000000, /* 3422 */
128'h1b0000000f00000003000000a0000000, /* 3423 */
128'h000063746e692d7570632c7663736972, /* 3424 */
128'h01000000b50000000400000003000000, /* 3425 */
128'h01000000bb0000000400000003000000, /* 3426 */
128'h01000000020000000200000002000000, /* 3427 */
128'h0030303030303030384079726f6d656d, /* 3428 */
128'h6f6d656d5b0000000700000003000000, /* 3429 */
128'h67000000100000000300000000007972, /* 3430 */
128'h00000008000000000000008000000000, /* 3431 */
128'h0300000000636f730100000002000000, /* 3432 */
128'h03000000020000000000000004000000, /* 3433 */
128'h03000000020000000f00000004000000, /* 3434 */
128'h616972612c6874651b0000001f000000, /* 3435 */
128'h706d697300636f732d657261622d656e, /* 3436 */
128'h000000000300000000007375622d656c, /* 3437 */
128'h303240746e696c6301000000c3000000, /* 3438 */
128'h0d000000030000000000003030303030, /* 3439 */
128'h30746e696c632c76637369721b000000, /* 3440 */
128'hca000000100000000300000000000000, /* 3441 */
128'h07000000010000000300000001000000, /* 3442 */
128'h00000000670000001000000003000000, /* 3443 */
128'h0300000000000c000000000000000002, /* 3444 */
128'h006c6f72746e6f63de00000008000000, /* 3445 */
128'h7075727265746e690100000002000000, /* 3446 */
128'h3030634072656c6c6f72746e6f632d74, /* 3447 */
128'h04000000030000000000000030303030, /* 3448 */
128'h04000000030000000000000000000000, /* 3449 */
128'h0c00000003000000010000008f000000, /* 3450 */
128'h003063696c702c76637369721b000000, /* 3451 */
128'h03000000a00000000000000003000000, /* 3452 */
128'h0b00000001000000ca00000010000000, /* 3453 */
128'h10000000030000000900000001000000, /* 3454 */
128'h000000000000000c0000000067000000, /* 3455 */
128'he8000000040000000300000000000004, /* 3456 */
128'hfb000000040000000300000007000000, /* 3457 */
128'hb5000000040000000300000003000000, /* 3458 */
128'hbb000000040000000300000002000000, /* 3459 */
128'h75626564010000000200000002000000, /* 3460 */
128'h0000304072656c6c6f72746e6f632d67, /* 3461 */
128'h637369721b0000001000000003000000, /* 3462 */
128'h03000000003331302d67756265642c76, /* 3463 */
128'hffff000001000000ca00000008000000, /* 3464 */
128'h00000000670000001000000003000000, /* 3465 */
128'h03000000001000000000000000000000, /* 3466 */
128'h006c6f72746e6f63de00000008000000, /* 3467 */
128'h30313440747261750100000002000000, /* 3468 */
128'h08000000030000000000003030303030, /* 3469 */
128'h03000000003035373631736e1b000000, /* 3470 */
128'h00000041000000006700000010000000, /* 3471 */
128'h04000000030000000010000000000000, /* 3472 */
128'h040000000300000080f0fa024b000000, /* 3473 */
128'h040000000300000000c2010006010000, /* 3474 */
128'h04000000030000000200000014010000, /* 3475 */
128'h04000000030000000100000025010000, /* 3476 */
128'h04000000030000000200000030010000, /* 3477 */
128'h0100000002000000040000003a010000, /* 3478 */
128'h3030323440636d6d2d63736972776f6c, /* 3479 */
128'h10000000030000000000000030303030, /* 3480 */
128'h00000000000000420000000067000000, /* 3481 */
128'h14010000040000000300000000000100, /* 3482 */
128'h25010000040000000300000002000000, /* 3483 */
128'h1b0000000c0000000300000002000000, /* 3484 */
128'h0200000000636d6d2d63736972776f6c, /* 3485 */
128'h406874652d63736972776f6c01000000, /* 3486 */
128'h03000000000000003030303030303334, /* 3487 */
128'h2d63736972776f6c1b0000000c000000, /* 3488 */
128'h5b000000080000000300000000687465, /* 3489 */
128'h0400000003000000006b726f7774656e, /* 3490 */
128'h04000000030000000200000014010000, /* 3491 */
128'h06000000030000000300000025010000, /* 3492 */
128'h0300000000007fe3023e180047010000, /* 3493 */
128'h00000043000000006700000010000000, /* 3494 */
128'h01000000020000000080000000000000, /* 3495 */
128'h303434406f6970672d63736972776f6c, /* 3496 */
128'h0d000000030000000000003030303030, /* 3497 */
128'h6f6970672d63736972776f6c1b000000, /* 3498 */
128'h67000000100000000300000000000000, /* 3499 */
128'h00100000000000000000004400000000, /* 3500 */
128'h09000000020000000200000002000000, /* 3501 */
128'h2300736c6c65632d7373657264646123, /* 3502 */
128'h61706d6f6300736c6c65632d657a6973, /* 3503 */
128'h6f647473006c65646f6d00656c626974, /* 3504 */
128'h65736162656d697400687461702d7475, /* 3505 */
128'h6b636f6c630079636e6575716572662d, /* 3506 */
128'h63697665640079636e6575716572662d, /* 3507 */
128'h75746174730067657200657079745f65, /* 3508 */
128'h2d756d6d006173692c76637369720073, /* 3509 */
128'h230074696c70732d626c740065707974, /* 3510 */
128'h00736c6c65632d747075727265746e69, /* 3511 */
128'h6f72746e6f632d747075727265746e69, /* 3512 */
128'h646e6168702c78756e696c0072656c6c, /* 3513 */
128'h727265746e69007365676e617200656c, /* 3514 */
128'h6572006465646e657478652d73747075, /* 3515 */
128'h616d2c76637369720073656d616e2d67, /* 3516 */
128'h766373697200797469726f6972702d78, /* 3517 */
128'h70732d746e6572727563007665646e2c, /* 3518 */
128'h61702d747075727265746e6900646565, /* 3519 */
128'h0073747075727265746e6900746e6572, /* 3520 */
128'h6f692d6765720074666968732d676572, /* 3521 */
128'h63616d2d6c61636f6c0068746469772d, /* 3522 */
128'h0000000000000000737365726464612d, /* 3523 */
128'h0000000000203a642520656369766544, /* 3524 */
128'h00203a6425206563697665642073250a, /* 3525 */
128'h00000000203a6425206563697665440a, /* 3526 */
128'h000a656369766564206e776f6e6b6e75, /* 3527 */
128'h00000a2973252c73252870756b6f6f6c, /* 3528 */
128'h7265206c616e7265746e692070636864, /* 3529 */
128'h00000000000000000a7025202c726f72, /* 3530 */
128'h5145525f5043484420676e69646e6553, /* 3531 */
128'h4b434120504348440000000a54534555, /* 3532 */
128'h696c432050434844000000000000000a, /* 3533 */
128'h203a7373657264644120504920746e65, /* 3534 */
128'h0000000a64252e64252e64252e642520, /* 3535 */
128'h73657264644120504920726576726553, /* 3536 */
128'h0a64252e64252e64252e642520203a73, /* 3537 */
128'h6120726574756f520000000000000000, /* 3538 */
128'h252e64252e642520203a737365726464, /* 3539 */
128'h6b73616d2074654e0000000a64252e64, /* 3540 */
128'h64252e642520203a7373657264646120, /* 3541 */
128'h697420657361654c000a64252e64252e, /* 3542 */
128'h7364253a6d64253a686425203d20656d, /* 3543 */
128'h3d206e69616d6f44000000000000000a, /* 3544 */
128'h4820746e65696c4300000a2273252220, /* 3545 */
128'h000a22732522203d20656d616e74736f, /* 3546 */
128'h000000000a44455050494b53204b4341, /* 3547 */
128'h000000000000000a4b414e2050434844, /* 3548 */
128'h73657264646120646574736575716552, /* 3549 */
128'h0000000000000a646573756665722073, /* 3550 */
128'h000000000000000a732520726f727245, /* 3551 */
128'h6e6f6974706f2064656c646e61686e75, /* 3552 */
128'h656c646e61686e55000000000a642520, /* 3553 */
128'h64252065646f63706f20504348442064, /* 3554 */
128'h20676e69646e6553000000000000000a, /* 3555 */
128'h000a595245564f435349445f50434844, /* 3556 */
128'h00000000000a29732528726f72726570, /* 3557 */
128'h3a2043414d2073250000000030687465, /* 3558 */
128'h3a583230253a583230253a5832302520, /* 3559 */
128'h000a583230253a583230253a58323025, /* 3560 */
128'h484420646e65732074276e646c756f43, /* 3561 */
128'h206e6f20595245564f43534944205043, /* 3562 */
128'h00000a7325203a732520656369766564, /* 3563 */
128'h5043484420726f6620676e6974696157, /* 3564 */
128'h2020202020202020000a524546464f5f, /* 3565 */
128'h00000000000063250000000000000020, /* 3566 */
128'h0000005832302520000000000000002e, /* 3567 */
128'h00000000732573250000000000000a0a, /* 3568 */
128'h00000000007325203a646c697542202c, /* 3569 */
128'h73257a4820756c250000000000007325, /* 3570 */
128'h0000000000756c250000000000000000, /* 3571 */
128'h0073257a4863252000000000646c252e, /* 3572 */
128'h00000000007325736574794220756c25, /* 3573 */
128'h00003a786c3830250073254269632520, /* 3574 */
128'h000a73252020202000786c6c2a302520, /* 3575 */
128'h000000203a5d64255b6e6f6974636553, /* 3576 */
128'h727265207974696e6173207264646170, /* 3577 */
128'h2c7825286e666c6500000a702520726f, /* 3578 */
128'h000000000a3b29782578302c78257830, /* 3579 */
128'h782578302c302c7825287465736d656d, /* 3580 */
128'h464f5f4f4c43414d00000000000a3b29, /* 3581 */
128'h464f5f494843414d0000000054455346, /* 3582 */
128'h46464f5f524c50540000000054455346, /* 3583 */
128'h46464f5f534346540000000000544553, /* 3584 */
128'h4c5254434f49444d0000000000544553, /* 3585 */
128'h46464f5f534346520054455346464f5f, /* 3586 */
128'h5346464f5f5253520000000000544553, /* 3587 */
128'h46464f5f444142520000000000005445, /* 3588 */
128'h46464f5f524c50520000000000544553, /* 3589 */
128'h000000003f3f3f3f0000000000544553, /* 3590 */
128'h000064252b54455346464f5f524c5052, /* 3591 */
128'h6f746f72502050490000000000000047, /* 3592 */
128'h00000000000000000a50495049203d20, /* 3593 */
128'h6f746f72502050490000000000000054, /* 3594 */
128'h6f746f7250205049000a504745203d20, /* 3595 */
128'h6165682074736574000a505550203d20, /* 3596 */
128'h6e6f6320747365740000000a3a726564, /* 3597 */
128'h6f746f7250205049000a3a73746e6574, /* 3598 */
128'h6f746f7250205049000a504449203d20, /* 3599 */
128'h6f746f725020504900000a5054203d20, /* 3600 */
128'h00000000000000000a50434344203d20, /* 3601 */
128'h6f746f72502050490000000000000036, /* 3602 */
128'h00000000000000000a50565352203d20, /* 3603 */
128'h000a455247203d206f746f7250205049, /* 3604 */
128'h000a505345203d206f746f7250205049, /* 3605 */
128'h00000a4841203d206f746f7250205049, /* 3606 */
128'h000a50544d203d206f746f7250205049, /* 3607 */
128'h5054454542203d206f746f7250205049, /* 3608 */
128'h6f746f72502050490000000000000a48, /* 3609 */
128'h000000000000000a5041434e45203d20, /* 3610 */
128'h6f746f7250205049000000000000004d, /* 3611 */
128'h00000000000000000a504d4f43203d20, /* 3612 */
128'h0a50544353203d206f746f7250205049, /* 3613 */
128'h6f746f72502050490000000000000000, /* 3614 */
128'h00000000000a4554494c504455203d20, /* 3615 */
128'h0a534c504d203d206f746f7250205049, /* 3616 */
128'h6f746f72502050490000000000000000, /* 3617 */
128'h6f746f7270205049000a574152203d20, /* 3618 */
128'h2820646574726f707075736e75203d20, /* 3619 */
128'h79745f6f746f7270000000000a297825, /* 3620 */
128'h0000000000000a78257830203d206570, /* 3621 */
128'h727265746e692064656c646e61686e75, /* 3622 */
128'h414d2070757465530000000a21747075, /* 3623 */
128'h4d454f2049505351000a726464612043, /* 3624 */
128'h0000000000000a7825203d205d64255b, /* 3625 */
128'h00000a786c253a786c25203d2043414d, /* 3626 */
128'h3025203d20737365726464612043414d, /* 3627 */
128'h3230253a783230253a783230253a7832, /* 3628 */
128'h0000000a2e783230253a783230253a78, /* 3629 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 3630 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 3631 */
128'h66656463626139383736353433323130, /* 3632 */
128'h72776f6c2f6372730000000000000000, /* 3633 */
128'h00000000000000632e636d6d5f637369, /* 3634 */
128'h61625f6473203d3d20657361625f6473, /* 3635 */
128'h5f63736972776f6c00726464615f6573, /* 3636 */
128'h000a74756f656d6974207325203a6473, /* 3637 */
128'h616d202c6465766f6d65722064726143, /* 3638 */
128'h6425206f74206465676e616863206b73, /* 3639 */
128'h736e692064726143000000000000000a, /* 3640 */
128'h6e616863206b73616d202c6465747265, /* 3641 */
128'h0000000000000a6425206f7420646567, /* 3642 */
128'h25207461206465746165726320636d6d, /* 3643 */
128'h0000000a7825203d2074736f68202c78, /* 3644 */
128'h0000000000006f4e0000000000736559, /* 3645 */
128'h002020203a434d4d0000000052444420, /* 3646 */
128'h00000000000a7325203a656369766544, /* 3647 */
128'h3a4449207265727574636166756e614d, /* 3648 */
128'h0a7825203a4d454f000000000a782520, /* 3649 */
128'h6325203a656d614e0000000000000000, /* 3650 */
128'h0000000000000a206325632563256325, /* 3651 */
128'h00000a6425203a646565705320737542, /* 3652 */
128'h25203a79746963617061432068676948, /* 3653 */
128'h79746963617061430000000000000a73, /* 3654 */
128'h7464695720737542000000000000203a, /* 3655 */
128'h000000000a73257469622d6425203a68, /* 3656 */
128'h0000007825782520000000203a78250a, /* 3657 */
128'h00000000000064735f63736972776f6c, /* 3658 */
128'h0000000065646f6d206e776f6e6b6e55, /* 3659 */
128'h7830203a726f72724520737574617453, /* 3660 */
128'h2074756f656d69540000000a58383025, /* 3661 */
128'h616572206472616320676e6974696177, /* 3662 */
128'h6c69616620636d6d00000000000a7964, /* 3663 */
128'h6d6320706f747320646e6573206f7420, /* 3664 */
128'h6f6c62203a434d4d0000000000000a64, /* 3665 */
128'h20786c257830207265626d756e206b63, /* 3666 */
128'h6c2578302878616d2073646565637865, /* 3667 */
128'h203d3e20434d4d6500000000000a2978, /* 3668 */
128'h726f6620646572697571657220342e34, /* 3669 */
128'h642072657375206465636e61686e6520, /* 3670 */
128'h000000000000000a6165726120617461, /* 3671 */
128'h757320746f6e2073656f642064726143, /* 3672 */
128'h696e6f697469747261702074726f7070, /* 3673 */
128'h656f64206472614300000000000a676e, /* 3674 */
128'h20434820656e6966656420746f6e2073, /* 3675 */
128'h00000a657a69732070756f7267205057, /* 3676 */
128'h636e61686e6520617461642072657355, /* 3677 */
128'h5720434820746f6e2061657261206465, /* 3678 */
128'h696c6120657a69732070756f72672050, /* 3679 */
128'h72617020692550470000000a64656e67, /* 3680 */
128'h505720434820746f6e206e6f69746974, /* 3681 */
128'h67696c6120657a69732070756f726720, /* 3682 */
128'h656f642064726143000000000a64656e, /* 3683 */
128'h6e652074726f7070757320746f6e2073, /* 3684 */
128'h657475626972747461206465636e6168, /* 3685 */
128'h6e65206c61746f54000000000000000a, /* 3686 */
128'h6563786520657a6973206465636e6168, /* 3687 */
128'h20752528206d756d6978616d20736465, /* 3688 */
128'h656f64206472614300000a297525203e, /* 3689 */
128'h6f682074726f7070757320746f6e2073, /* 3690 */
128'h61702064656c6c6f72746e6f63207473, /* 3691 */
128'h6572206574697277206e6f6974697472, /* 3692 */
128'h6e6974746573207974696c696261696c, /* 3693 */
128'h726c61206472614300000000000a7367, /* 3694 */
128'h64656e6f697469747261702079646165, /* 3695 */
128'h206f6e203a434d4d000000000000000a, /* 3696 */
128'h0000000a746e65736572702064726163, /* 3697 */
128'h73657220746f6e206469642064726143, /* 3698 */
128'h20656761746c6f76206f7420646e6f70, /* 3699 */
128'h00000000000000000a217463656c6573, /* 3700 */
128'h7463656c6573206f7420656c62616e75, /* 3701 */
128'h00000000000000000a65646f6d206120, /* 3702 */
128'h646e756f66206473635f747865206f4e, /* 3703 */
128'h78363025206e614d0000000000000a21, /* 3704 */
128'h000000783430257834302520726e5320, /* 3705 */
128'h00000000632563256325632563256325, /* 3706 */
128'h6167656c20434d4d00000064252e6425, /* 3707 */
128'h636167654c2044530000000000007963, /* 3708 */
128'h6867694820434d4d0000000000000079, /* 3709 */
128'h0000297a484d36322820646565705320, /* 3710 */
128'h35282064656570532068676948204453, /* 3711 */
128'h6867694820434d4d000000297a484d30, /* 3712 */
128'h0000297a484d32352820646565705320, /* 3713 */
128'h7a484d32352820323552444420434d4d, /* 3714 */
128'h31524453205348550000000000000029, /* 3715 */
128'h00000000000000297a484d3532282032, /* 3716 */
128'h7a484d30352820353252445320534855, /* 3717 */
128'h35524453205348550000000000000029, /* 3718 */
128'h000000000000297a484d303031282030, /* 3719 */
128'h7a484d30352820303552444420534855, /* 3720 */
128'h31524453205348550000000000000029, /* 3721 */
128'h0000000000297a484d38303228203430, /* 3722 */
128'h0000297a484d30303228203030325348, /* 3723 */
128'h6f6e2064252065636976654420434d4d, /* 3724 */
128'h00000000000000000a646e756f662074, /* 3725 */
128'h000000000000445300000000434d4d65, /* 3726 */
128'h000000297325282000006425203a7325, /* 3727 */
128'h6e656c20656c69460000000000636d6d, /* 3728 */
128'h000000000000000a6425203d20687467, /* 3729 */
128'h0a7325203d202964252c70252835646d, /* 3730 */
128'h666c652064616f6c0000000000000000, /* 3731 */
128'h000a79726f6d656d20524444206f7420, /* 3732 */
128'h2064656c696166206461657220666c65, /* 3733 */
128'h000000646c252065646f632068746977, /* 3734 */
128'h6f6f7420687461702074736575716552, /* 3735 */
128'h00000000000a646c25202e676e6f6c20, /* 3736 */
128'h732522203a717277000000000000002f, /* 3737 */
128'h0a64253d657a69736b636f6c62202c22, /* 3738 */
128'h20657669656365520000000000000000, /* 3739 */
128'h0000000000000a2e646e6520656c6966, /* 3740 */
128'h656c6c6163207172775f656c646e6168, /* 3741 */
128'h206c6167656c6c4900000000000a2e64, /* 3742 */
128'h0a2e6e6f6974617265706f2050544654, /* 3743 */
128'h37363534333231300000000000000000, /* 3744 */
128'h00000000000000004645444342413938, /* 3745 */
128'h25203d206465726975716572206e656c, /* 3746 */
128'h000a7825203d206c6175746361202c58, /* 3747 */
128'h65687420746f6f42000000005c2d2f7c, /* 3748 */
128'h206d6172676f727020646564616f6c20, /* 3749 */
128'h2e2e2e70252073736572646461207461, /* 3750 */
128'h206f74206c696146000000000000000a, /* 3751 */
128'h2172657669726420445320746e756f6d, /* 3752 */
128'h6f6f622064616f4c000000000000000a, /* 3753 */
128'h726f6d656d206f746e69206e69622e74, /* 3754 */
128'h6e69622e746f6f620000000000000a79, /* 3755 */
128'h742064656c6961460000000000000000, /* 3756 */
128'h0000000a21746f6f62206e65706f206f, /* 3757 */
128'h69662065736f6c63206f74206c696166, /* 3758 */
128'h206f74206c696166000000000021656c, /* 3759 */
128'h00000000216b73696420746e756f6d75, /* 3760 */
128'h696620646573616220746f6f622d750a, /* 3761 */
128'h6c20746f6f6220656761747320747372, /* 3762 */
128'h6f6974726573736100000a726564616f, /* 3763 */
128'h6c6966202c64656c696166207325206e, /* 3764 */
128'h66202c642520656e696c202c73252065, /* 3765 */
128'h00000000000a7325206e6f6974636e75, /* 3766 */
128'h3d212078257830203a4552554c494146, /* 3767 */
128'h2074657366666f207461207825783020, /* 3768 */
128'h2c7025203d20317000000a2e78257830, /* 3769 */
128'h000000000000000a7025203d20327020, /* 3770 */
128'h00000000002020202020202020202020, /* 3771 */
128'h00000000000808080808080808080808, /* 3772 */
128'h000000000000752520676e6974746573, /* 3773 */
128'h000000000000752520676e6974736574, /* 3774 */
128'h6c626973736f70203a4552554c494146, /* 3775 */
128'h696c2073736572646461206461622065, /* 3776 */
128'h2578302074657366666f20746120656e, /* 3777 */
128'h676e697070696b5300000000000a2e78, /* 3778 */
128'h2e2e2e74736574207478656e206f7420, /* 3779 */
128'h0808080808080808000000000000000a, /* 3780 */
128'h08082020202020202020202020080808, /* 3781 */
128'h00000000000000080808080808080808, /* 3782 */
128'h6e617220747365740000000000082008, /* 3783 */
128'h7830206f742070257830207369206567, /* 3784 */
128'h00752520706f6f4c00000000000a7025, /* 3785 */
128'h0000000000000a3a000000000075252f, /* 3786 */
128'h00000073736572646441206b63757453, /* 3787 */
128'h00000000000a6b6f0000203a73252020, /* 3788 */
128'h656d20657261420a00000a2e656e6f44, /* 3789 */
128'h00000a74736574204d415244206c6174, /* 3790 */
128'h7025203d2029286e69616d5f6d617264, /* 3791 */
128'h287073206d617264000000000000000a, /* 3792 */
128'h65747365746d656d000a7025203d2029, /* 3793 */
128'h20302e332e34206e6f69737265762072, /* 3794 */
128'h000000000000000a297469622d642528, /* 3795 */
128'h30322029432820746867697279706f43, /* 3796 */
128'h2073656c7261684320323130322d3130, /* 3797 */
128'h000000000000000a2e6e6f62617a6143, /* 3798 */
128'h74207265646e75206465736e6563694c, /* 3799 */
128'h50206c6172656e654720554e47206568, /* 3800 */
128'h65762065736e6563694c2063696c6275, /* 3801 */
128'h0a2e29796c6e6f282032206e6f697372, /* 3802 */
128'h5f676e696b726f770000000000000000, /* 3803 */
128'h20646c25202c424b6425203d20746573, /* 3804 */
128'h6c25202c736e6f697463757274736e69, /* 3805 */
128'h203d20495043202c73656c6379632064, /* 3806 */
128'h00000000000000000a646c252e646c25, /* 3807 */
128'h524444206f7420495053512064616f6c, /* 3808 */
128'h00000000000000000a79726f6d656d20, /* 3809 */
128'h20524444206f7420464c452064616f6c, /* 3810 */
128'h6f57206f6c6c6548000a79726f6d656d, /* 3811 */
128'h205d64255b70777300000a0d21646c72, /* 3812 */
128'h73206863746977530000000a5825203d, /* 3813 */
128'h000a58252c5825203d20676e69747465, /* 3814 */
128'h5825203d2064656573206d6f646e6152, /* 3815 */
128'h0a746f6f62204453000000000000000a, /* 3816 */
128'h6f6f6220495053510000000000000000, /* 3817 */
128'h736574204d4152440000000000000a74, /* 3818 */
128'h6f6f6220505446540000000000000a74, /* 3819 */
128'h65742065686361430000000000000a74, /* 3820 */
128'h00000a0d7061727400000000000a7473, /* 3821 */
128'h00000002464c457fcccccccccccccccd, /* 3822 */
128'h1032547698badcfeefcdab8967452301, /* 3823 */
128'h5851f42d4c957f2d1000000020000000, /* 3824 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 3825 */
128'h000000004503e0000000000045030000, /* 3826 */
128'h000000004503c0000000000045040000, /* 3827 */
128'h000002000000019d0000000045038000, /* 3828 */
128'h00000000cc33aa550000000084000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00004b4d47545045000000030f060301, /* 3840 */
128'h000000004300000000000000004b4d47, /* 3841 */
128'h00000000ffffffff0000000000000000, /* 3842 */
128'h0000646d635f6473000000000c000000, /* 3843 */
128'h00000000ffffffff00006772615f6473, /* 3844 */
128'h000000002f7c5c2d0000000087fee748, /* 3845 */
128'hffffffff000000060000000087fee900, /* 3846 */
128'h0000000087fe709c0000000000000000, /* 3847 */
128'h0000000000000000000000000000005e, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule


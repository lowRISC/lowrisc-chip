`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RfRAPnyT7kS4fe+DSlNjyfm+lxLWmnOc/+s3ca7Kfsg+t2gE4bq+JaYlQDM990HI9wpRT6ORcXMv
m4QvOTEkqraxDauZ6pEjlFZLAWkBn2RD+Y68tSsj8j+r9cdBuZSKQmCD186SeiHn2n/c71cVvhCz
0+vLYZQMFF1s/V1Mqav7bLWzehoGtbAibBjUpIBNMbAthrhfl21w7DJpAcOPd7pEWw0kgLDBtwQZ
738d/VdIVwDOei1ulmKD4znQz9KnE9bYEWc8v0PLLXNN/Za78isNEtPu5LwL5DJtzgNek13z+oRo
FqwA7vMJnxzhP1NmKgpYplaOlgT7AWj2bZ6nKg==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
qWnWJAQ7xuikC20h3BRVNtsGWDO+zlQHYMOjScKd9eAv48xkJH21xvDNBycUEAyvVxRnhkXvXFk/
09U8wWAPNQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MpyauYkejEmNftb97dhw4aGFKV9W4EQMtkPpjhhdHJjGjhUEzCXiw5ZlpzxTU6scCIN9zO5tHEUl
jsVxjJaMAyILTQiz/S+DiliunK+fX79en2xXjX7WszdDBp37sgmyECfcOtBab+3pixTC76qkAn4B
RLXQUYa4FrFmXDnqZb0=

`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eakjADqkxZxvMiiOcYpslfNYhD4gQfH863GOmMA+/yi8fcE6aKcfFP+cdZ3PCgzFTPxKXh4Xo0qO
vSYqymGdYR3PF8no5g5hqatU3ArRfpWMXFJqO+qjJ5xFJRf9uzFFcgDQfAoqOamQOLuJFsDGHk7O
e0FQ9P57AOaCvjh59Bg=

`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dm1AXsH0tpajjYg92+oFVNb8hBuDxolZQNjMj3a8MeCl9VZjJT1doOVBIKT1t5cxrCT4QSXto/1z
Z0f6CGXGy4s1T4HXz8JVS/rP452MrEcsA3YVCdTBrlNfqvAwJzSyjtZgev8BulEbPGEZMo9Yji1W
HRCuRPSLKJbk4L2WumI2956bs1ZNwP2a+7SEHSHf9VrOMhX5KdVbmdS9nSbnoP2DLkNiqoubJJ5S
+An0XyzEm4Rl8zztbfj4Rpyeac6y3QDoMv0na89VoQM0raK7H0Z5iM4s+MUaLs8yGptPFO4A09T0
/skipuXt326AVG+m8ZWF7giIMTBy4ldsCghNsg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135632)
`pragma protect data_block
C22JCRackNK2Z70cE7Q5xToQr1s946xfcdZJ/3lSt7y2OTtgAgeP9tAAxZxvyL6B9AbfUjExvytc
SxyJcDZqJ84udOSK6G6rv/V8hS8RbIMJr7wl7ht9Celv/GzJo3ox7ZgY2QL2ddhMIh2xr3OEBr9I
RfxmmtZ2MsQiA6SbZ/I5+09Qq4DD/6za7kBzC7xoxqy15RJGjFEQaRPT9lOgh13U/YBYtevzE5gW
PVfv7a6IOmYBmIu4a3rWEe6IaA+J9DUO6pW7HMncoWSQatgq3a5XbyaiQmrryxJIRFLXa1NwPOen
mdag5bycDZMp63Q7oXtVbR5wOPC3i0NcVVYjwMnDo15ZAK/ECOORsoawczj2OAa6ZQaJT+UcTaws
5i7+xr7m+ZoaFL3YDo4wcAuuf0CSITe6AJNdDIQDiu7YW/UIobpdNPfSvCrJQvvZBO7Q4dUTt71y
zDssA9fw3ldT6seT9wZzEn+ai1KnDXhAkDn/MFGqeLQSUeQNNZ7Dr+AOMde5Td4nOp4gITsQFbok
RKspI65HahSfL+GrRbOmKoUFM9hCwkhOoj0u+TVHkKD54G/Qy8OdBIZu3T+0CVxsMvm5ONwR0/DA
651w5YFDcU/msPqD+SR+hheWK3Ky+ycsN8P39zCjmSIm8Y1yelV95UfPVtNFuBMz5FubP10JK5e6
a2xdrAHHgVg0ZALhsEXTvdPscRV3zJKYEng4K3lwlm6EzoW78tW4Z6YCV3c8nAnqFMl2ZURy+LGh
uILsVL8T/eBSVoAn+uCONlpDwvOvI+I/N6Ych5XbWZ5L+NjnQsPLJ4sLx3ACLrM1la57rh3VQIHr
ERDEVKPGZ0RzcM4DI+/yGQIo+VO7u9fMfiIV3oIAbr3Ivn+0gDTyebQ03U3OGDjeKQg8lEIDxllG
RQzllaeNAORiLRphFhEuecTlj6U+gHKe275h1eYWUWDvkXzbFcTbZwcEcWJEw4FVpB490m272xGI
hJ6wbYu+nC+8WRMht7hhFmXAn0qSjFlspfddt9YhqFKPyBvmh3otR4sz4IPCYyNNRI7BP6gOgpcs
+sWut1rrft5MTFT+1cJZStZePYKz1Jxf29UyA/icfTZ27jxwa6SMfE0o+rjqFf9+f9IKvjxclX0D
8OE/e1VGQbB+3rGIm2nFlCw7Tu14ITf5g4fIK/ewGxsjdy8bnTuGYJ+gnAUAJs+6/vMFvbnXAAIG
BYITUYTA0+uh9lmIBW1qJuZcWpMvSDJTpNLZEHIa2M7pds70ugiJPQg+d+VuXq2+3WPBTdbIwhwl
9LhOZPiZ5ifFCWrhweQYAQ6GCS6187XFNJGWIJdzTDwRG1Uw2h1mxXDCn1UYdUNLPvEKfu7+JPc+
/fNrqrD6PICmAs9QEIoU+TKcUF20494nGPU/FkavXJPh0UKYAsBpTYu1h9fozI0QE9sBuCUgPNiT
9Mvr8jxZEts+Hv/7PBhBrsf+08sqcD9BL/jCzyYeKTGwT2FK+r8EMEjrK7yYkWKq9BiykDyZT4l2
Ltn/q8bQq0H3QN/sc8qjshXSN0USU+a9EpB3oKevj0JzmVRxa3SIlb+BVvJeGPF9IDJN9p4ln4mB
lvkbhOam2pADJuIfPJEy1I/120rYQtH4FuXeWIHyJIepn5u+dxYYj2DVyfT03QTDaHUKPdZqCC7F
6CXtkKmYfb1Gp/b9nYEptxJYyOA+PrATEBVC/r6qlxT8IHJGhB7CvdQX8hFteo24FoAnglcGiW+N
Pu2jmvVQUvMLXedhwyQ7NsrXRWTrCH9KbdSZzfrceclD7cx3ng+XRXD9uWGbccePRKeKfB1ZWWzm
Nsto3TV2Qq/ef0xHn98sKcT86SaURUPbMXmBmk6ZNlc+Rwa9LKu05bNome27a29omAYsDlzCWvnP
1mW7jquYIVbZw6/741PDI3AHbKlruh4kTtT1N97yeD+R0C3DQGACBSLmrUqinGa3l6cZNaOFA8uQ
0AdjPLQzvQfnkCk/Wj6x1oIFFxYZHwkJXswbaj3CUYuFM4WQbQUbhinlaBho69W4Ln3P+q7yKX+O
twBFqDXxzStv7oSbgGhFZiXmr/wFftiY1locZwdvrfqwjG6UJc7/zs28KSRhW4qJHVp/vg+sYt2D
Vm8HhVlJQQvKSM32/c+hK1L563RrykeqPmK/z8w/jdkZasPzUbKPNaDk7ri7mlpWAyBwS3+AqFuf
ypcTzCw0eFarisPbRrwv/xkUiUNngaZweapSVvUmYQWE9seN9rxVT/wolFQZIC0WWLonvKSAHht5
wEWTt6caUZOJsBsLjuJi0WarThxnQCZUwTFRsJp87aRMgbNNekQrAOum4BtohXSxQ+EtU2gPxAwK
RKXA30lZ9CygNOHUem+D0bQ8y5pA/l1O0e7WaxMHUpmBBaTa30AaJUSBtHo7oYNH2xuWd1tLKtnR
vv0EmkP9Hsb/NctOpBSP+r3IEyOAtH59skt6y+B9kZ0H8wxCaanFIEJNwsTLhpHGqeBn9Szar1Z5
aTjtpvRjfGC8Tz0lTD+zlvr2PvV2SHldvCZFFTvIfNxfop1CvMmELPSm+OMORaObEcM31OROJTWn
1iqtDX0pobLtbPcD19HSmLmShI6QlH9uklLLN/ztXuSAdVq6z1+eAFGoRhVezQL/nwSAidFVtYFp
C0xxMCRTXCjHKwnH0+JY2kuUHJAQ0jZ3D5fwKTWrvgLJLwYKYSdPNkZPjZq1ExCF36WlYyWJKebp
am4NjajD0ZIYPFYHBAe0F3a2nzluuTawFpKLQjR5UgMGEf9Jg/jQI0gHKx2QapmUUKSok7SSNGDf
5fEzLuO/WdOs+7EP7nluw5NziJXtq2u9y1GSf53nh/ebzzByKBBWnMfhxSqNy8AbP3Roq8FaVcLW
AjpG0XJWe+erK7gSQuXNzlkU6rh+qWkP+bJ3U+0JQeGeFKYb3pwWPc7jKLoWFxTSl4QdLT3Tg+f0
ilUzHsYR2RKxvz02e/rNIXQUmrIFW+Fj5Rd2gwPmHKsXCePXbWsuHLPuGGvWK067W0Kr5bk7tkcn
H5dprgESKXNoID85Qc/2/vqAGrU0lNtn2K6AR6fjLKW9HjEj0vZqvFZ3vy3bqSdHs0AfnpqiTI+D
o52n9+Ng1G1dQsLn40jypS4rErNKgFf09WoUcVX/2R0a8C6cOR28+qAviOxJ8PZ5FfpKSl1JerKe
F/j584RCqSumtHJOPA6QzkLXtk/6yX9AI5zgsO5+HtJHy7XjBEoOOfJjglkJFlMuPKWebuOFf5xW
7X7+Fjc0yVkUDoZwAUReCFL+w1+/rT+BvXineO6SZ/zuMl+JAwD4Z6i5Z3r1W8/uk64Yi5EsFro2
A9k0fRGG31g4N6/e0GMYERyEJHOHSYNqypwMqGNpsDqQ6zT/IZ/U1+16SVRC2CoVdiV9IipH48lu
di4QLGUc6+vXusReO5/nHUvuE28jDbxZ/IOm5H35S7YSUVobcqCXO+Rool5YaDR+7zHYpPH3HQ3f
jWzHhpCTeK6Swj+/jYfuxUn18OmszRX+BsOf4mDFOYBSxUyX8peYwj3DFHnb7T2ga/aj7UTI0MOf
MQl6QZtHiUHyuYn/jYXtBOOihdq6foeytUOlbM6ZTzj2tpIW5X0QKEofF4I98ipP5k+MXr2G0aI5
W7X7KTCQ8CiMXQAGIgSz4wcGiuvR3cODLHWGERuhoD86u6bNNP4Su5fBU0EANjEfkzh95usMbYOO
h37lfSnl4e12Qb+2yZWMZ58cCkiPhYwqj2FK0aRTTsXZVZqrV/Y/5mQuAkhN3C2gs8x0yS61jCO7
H1+U6t8p3FE0oI49XtC3Hbu+CF9OkSXiVINVCZZ/NVd14/ZMEL6UEZkBu9yf4NYEh0cq5fOHjWiF
DUsCiSAzXC5p39xH3httCCDNnUD/uqj2lRA2gzUxpeBTxt5YPCTtgfDl7RzEeoafSS8uln0SYA/p
IDJwavxfJe0Pe45HLminU/25KF2I3g5Oz+SC3XD/rWL3+Y1XVm88UnC6vizvy57vaNHdpUGbX2uU
q8WWCUDEpuEaOAazJdza9IzLczh5wZB3+kcudX/E3MSkXGPw1LvSmLF/zIG+h12Me/S3QF5RE4/s
fnGRcO1M8IikszJVndnNZYcEnctn7N14M//IZDQLP7MwkkaPUQJKgSHrttHbcW/nJiuOs1Lt+LKt
zurNuzqVxfwm7+HWFRA/B4SGFdE2C0FJ9KbxRfli7rtBb7RXTmW0Kmhykdfuy2LrMBtJlUS9rnc/
iUAXdC7c5RlrkSoGQo5qZz0NTNJ2mj52fhdqI/ZdEUxqYsh6osLGPt9uX0ADEValAktlxKgToe6d
/SY5NbWF+r0tuseCTGRkQqILewRF/CXh265ay3qCn58UuxFrtej08CI9i8K5rGf4W2iGUbGOx6lr
eiI/xXCVHEqOCgY0WIAWDnBjJheTRSIgJ0I/UO/JzLrxM9biXh0DayIF0fNqbFdSG0Y8H3BskFCT
rUhSMjfAuZrfHcFgLhA7TG1D6kXMnubeq6HYAPvJv7bUWjBNT6FoHjPKn71xqe8iSXEW6Vbajbnu
gCclxYxSxUcFgTbeKLq2K8pIcrBtzAwNUs7WYlM0UeigjAXeILKKBHGtOfryktzxYnTlZRRtndgG
CCEqUQav0418rCfauOgFVg+2NMwo2mHLc9pjODorWBdMT4C7wPg6fABcDFTMtCV3Wn7t+aUerHia
lqTnYDMLr9O97WoMaq0aGxHJ12Rz1nSsNkYQ2Eqo6OojyfIrZ6RmTXDfMgp2aQ25NGrPeLcmnHQC
zqCHoLKmmcXoWPjbQxhJ7Cgq1bn+g37NqgDfqaCnK8H/mFt6DrWjMYDH6e5vHUuXtJDSojl6MtJ0
pwNnaAwcInwOPiMxU+M7ZvdzYKIfaw63eY/iZBZTtFwz/q6/qdHUSLPNDyQ50zVsVStKq0uUFhIU
CBSOnm4cSvNglk9Zv2oegEoiNOUv8A67ke3W7QrGS3MKAxO28xH/dJOd9iSTMOhFTBMYwN/tXoXk
iRNE9PgmJRCdYd0KCAXTqKBXiZXb45jyoBPJbLax9vSxpM5CmfYMN1OMymuBLLauLYNnl4BqlIdi
YSBhZHo+Tzm8zr6nEMbOfNQkyT8KgRumY8jNyKFUmRz8c1ugIkEceQary+b0dPZxVcGlw2poQ2eR
k9pJvtitddlvbT04L400cQc5nkgzuJwFHJMfbZRjZ+IE8uO/zSTfNF+v03fGX0vMmrF61lpG5d7m
hFZZqmOQFUrO+ds+rxIz5CUpy8uIRhfGJSqMKnyjOk2L7MO5Wnh6S6jQqp8NYVpyexwRUtYSzzOK
OJ3w4fdUjgjiFZrXXvmQl7hdNq6B+wDvJj6ACnUI+oR7q1C8wLtx1HPQcoSGuJ94vS0TNCY7EYFE
nN922GcELcJjRDokLkfKLammN9mzKXiEjIPsL/fasoVuwy5DJA9PuWPu3IVwPmD6JPQ6q9Q6Td8u
UtlJh/Udpc/Vzwb9aP5za6nP96t0XbrfR4vQIJMEvkWqcch/WyZ9bU5trdtf3S5FqWheU6Hs5D/6
JF3DOwbKEidV4kRU6Hnj4KQ6YKA0wMnQYSikMc2TBG5URYscf1vXrsclliy7nQx5rc9XZD8lFJ+k
3GuvhQuW9yXp3WMZjaEuTv0HUpE/tb5zWM9e5i9FmbNs9CdGNJE3bz/AVW9TisEmj5x4WJnBI6lD
Qt12QyBKAv1F+sFVFw/VYXPCrEYHiA/VMzQsffvERmqr+aIM2ymhlgGTng2bL8T9ZoKZtDJKnApp
AOdQNk82As9KrpQy2rfs/8V84qdSwkCoyhYEksRsNPApBj1TyKOMKcCJ546aXXZh6QoIAMBvw+tD
0n8Hgo34gJ8pFfS4hOvtBngiRWbkGWfkyX6ujLTpKxEPtv8c0LpaO+Vi4Ijyuo+DZt9dJI/MA0qP
q/JP4qy1MjAyfKoJMfnUUgs3FKpXHPe2eqrlOvJgltJbXMrrX2BAxK4k5sz4P3phZFTAPQ0ilvaC
qKmSE9pOKpBcaKnR1MWSoZ5miNnNPFA+dRm+h6rUdA5noBjtq6fsXO9yu4myEhEHoTQVuw9j8VZQ
rr5YjAI4HqB7GKmAjvfFRyC6deWWEwFbQmYsHqz/0ZSjBPOIKe/UxFXpxq9r8FhYJfu11IQSRVE0
E9XcPx3IYlHaxugywd2iKcBkUEyZdR822feWYMcOY2zscKktDWagfqiwVNIwiyd6uXGM2oE3DwBE
XgG8KX6Fprb0dFWW4IWLpV1+ektYA8csbX+yDIj3gEWWOZ7s6truOYkrdC1RgbH1fwQ/NbIbqT5X
3Xw89co9vRebh8PrEJdyL67TPb66JbOW03JMQmGcYICPIEvBX+x1JNh1FOGRqPf5fIwdthu0IvjM
hK6ecP8U1ZlLz2PjIrpRAYXZl9f50vCHQ81MTmz5dqU6ZpB9eor4mOFJvwlT/O8Di8rDrKjLoqlt
usOchCvisxcmDejNVjuEpMjplF4zFrz6Qg3vjRdRDHk8w32GARC8We4f+Cu9DiiNljpszA828Kxa
2AOPHKh07JO3T97P6C9AusCONOV8jKTMLgQ/kNILzd/3YMZulavZLttC6A3CZu+gxHSC75PdVGBu
c5IVWVSPhcy4y80mIwwvhE8gSY2yfhGfOo6w/1GUfFNRPG07xiOcedZfdqbDDrR6D2W92JlF0EG8
gQkkso4dm9g4TzwXqhsoUwi/D20+LNvxhiADD/cA4V8hqv5XqYtrDm+rxvNDTUAeLPS8e0plZz5m
CS4g2xntCT34M/F2YDL6n197LAER8OC4LVFLNH32+UKDAp0ASx8UC4utvBRnoiL1pm3nhTYvaT8l
8zPOw1PkK52jADa5BTH7BuOkvlUT8fcL7idhcqxU33vptVTja2QBp2F/KHJO7zY1aVb4at6jMm/N
88G9/Yhwu6zHBLw/1MSdMtGPfkyHS4qfhQJTEqRZGLzWfUSxZCM/WGrgWPMpCYLImTG+iS037rR+
oEPBX41nc4mvnurMm58Up7I0ejmXWqjTW9nJtFv5t2ZDkYBIPEzOwetXwWmwEADWF+NxzXrBXeLa
y2Q8vhAIhfxSYf49S7NMLulo7PTGUNrlIiAVotc3enWad7RAUlDYzTAHv/mMed7n11waznlGmlDB
qBgXxl/xo7IjNU76rUTwIeLF9B6rsaeBmzHY1yaHmniDS7fWNm39tmBX/CKHCGwtlCwRsH0rlDbp
xINzlsiZPY1ZoIytpiWx60+/KTVB/B4k5oXcCztdAAGdwwIQRHapQW0N/QCOfITYWwl+sxQsn3J+
cO+nRlbjH2btWmgevugNRD+ZwNFHM/dbxCCtsVdwE8r6f7YVKzBm9qAoLBfJJ7P1CwR1cTtcgg7L
aqX+nmh0hpB+AJiqa6c6wIibnLVdx7VyNR9CbU8U4Iyq+CpNI1iWHjnQaZhF0XjCffPKqK2V2Q8i
kZSr4v0jW5f8tMpm6AZWMLehCTs+hox78IQpd0DuTji3mcatKvdbSz5ietr6nQy+h/8iA5k2OQxs
nocpeh5pNoMo9Z+zUKUusWnHcO2CwPWFtcW29cYHaiDYfZkX4G5Ok1Wy63MBLZ/yItO4GCwkVQE6
oh/S0awU+MV9CP6AX8RFplp8zfgNmK73yIeTrX1NIUzzT6QQeLva56TdyYTaiKRWfNA+nqjaYCJa
LbyC/SaScpono7iDeWOOOnVj1AkZHcQ5fmwwpgiS2C1yOYQ7kC7EK/7+hFPH+G9gqc6SDy6Klxso
fskzXojb5gQDKB+rYF3jq9ultpaB/sR5kgru2SJ19HQ19IgXTgOA0k84rVFSpNBmX5F3Z/zZ6kkx
nK03i2/LXaRu4oOsmBrb7599onouuRSoWKs98vz/tdWo7oMJCjQkagjkXl6oc3k74IIXKI/3jc0a
5yhKE/gXqw0WT4nDaz0uaFPI6McA2fr3bRs+t9oH1b0pEmk1hyKKuEfYeWZGEnOXxzVqVm8h/MAF
FvvgKvgXD5JgkPTLJuWdfCDHr9GHwt6XNQVhjm+b45GpOrn81Kd2u2mKLeR3zD0A3jd91oJBoByp
ckemP/O9qZmpMtgEizhKiOwvg64sfWkZ6H9KKWVAnNTwk+FIaAGU+28VQ3ntDWJymtO3U/Rh/sJS
gAoCzLCRyHJ63iyoOMdAeYSsZTy+yp32Zrmm0OHB3pl2lZjvV82fWIIIZStccu7HcQvZ+neYvt3u
rJ6UnA4uiJENkSBTLzu+frewLB0DkPq5a1EaoEfMm/ZWcC4bog1vWxGXC3YZ2ijGpvDJeemCvc7M
kLDgFAwc37/LWJx+gWRBEJMmnX+uQARVO5t8tikZF1armQyyWpvSNJR5OxBQKxRyxoCyP4akreEU
ceE6HJlXjdqbzq9SoJq3rxMm1IiOuzaBKCwUZsL4EEE5oiYPzwnyok6P2S9xta+5T8v/4vvVHcTg
oYFMLGaM3Sxvp8SU7fy6ydsY0fmWDcu2m7hEMFSA6f0NyYam/t0ViTmwZqJ8D18nrVWsKlO995wo
RT4SWY4wzka4NB/yNd0juB0WVsTNHzfc4O8MqyWR6phLJWTGd2HtaNnKIHAPn3nb8MR5tULHfE3F
VW9pPA6mn6mG3g7C12v66PKyDvaDrJbDGCjAIKbeIHynfQN4OhOYzzrirwvczxRT/agETdmnDVjF
NqIwiU5gEoAyB6aIHmFZkkZumRu/ZI9G/wiIy0sXjRxnp+uStY7soBwr6Ws9Q4k9A1Bq5VbVwsI0
UsEqF9uFBAo+bXaDJ+bY0qzEGKhnph5t+bICqlFCYKuY1DXCezt0RVmX1ZnwDSvsNldmtdVxRQ/q
fvhspi1ZXg/5rPSDpKo7qb9nQuE+XutC+8aIcpeM9Wia7z4vmMWWL7VcmiE1PrDsPB0aikIi4THT
fQV4GXHTxO5ycvW+AnU7QfNIweKS0mbbqGXV34WsMmPLodIlcQO6AszzhUZMl+av3fiNl4GmGMbX
hPPwl7cKOZYBMA/WX1fWt9jccGqJ1fmbNSaaqSFE+WSHxrHtTAw6CriVxZxlWPENY2QjEuXCjwPk
g9M2/Ruti8KemDCfcY0/Xv/nZ3SFdDAqDq8kZ2fpKNSOvCi2MOvDO/EOU3X7R0PGofs10dqyh+gZ
/0yLgfE5YXlIs4iSLnZZwugHs+yO95E5H3B88QWpw0VS0oRdIBV+EjclRXIEnBA82rhsX+Ms7VqP
+Iz5gJnGfz5WKTkgqwixUdYaC3Hr1WWNRSadi86mSVFQTeWkUznA0o52eFQIR8gb9tve9nHECuMZ
hsnk7UPnIPLKfXgnNGlI/gLQQyrWE9PFwfwgnIlSjcWHNyPXm2JtBDhdOEZmUXyBSjf979QNpiGD
KQxQKDqLFviJKJY+Pr9LjYM01j9FRQjI0NfKCq6kcpEYvuxx1iFALqC3c80+SVodNrnN/GqFk0Wz
o5j68382bouBEuGY9np0RDjiFuK+x2KY1O/J2veVkPdZEaB/170NhmnPsDwwWSUJKfjlLpRYNtvM
BKcB+y7RM3yUgkMWIh+jIk2j21lqR+pBIldNmo4Q1xl7/DV5PsykRA08+0TKRE2jskur32axA1DU
AgwUh0odKmCIAaf3+iPjqdhH8gaGcyGNZtFMTk0Q2ng8d/gf/D6Spb/xMkjn2CJRJhm7iLYrkqPd
t1CoV5vDcM7li9q9+e1oKdI8vrRSGJfRSA33mh4m8/tV8Rv8kegTn07I12zTa74SrPwGDzGcSKot
zNQCuHDkE7Am0SuGkSaFYinFmlc0jKHyfP2QfjXNKqbp01BrVhHPHxaOhd+f5sW9RQkJfjD0YhEB
2iDeIfPA/WkzOu9y09F3JA6mSBSH1HyZ01FgGxRVtS2gSEnS8Ic1fb0SajoPQqHfairla1vednAY
YsjplA8hjH4LL/GZ99wQS6RqJn8GpHexTsgT4d2n1VEnsKZYtiiyi+V4lSGIVH5NsqJvsfvxHh7S
57xhBiGMY/oRBxROUXIslNyIFePgKx6oPU5Jlsnbb0zgmepBxds/nkIlg0rRdILPKA8ScTTKu8TG
fbd2HvF4MHvNwnps5Iyep86KnFyFLog/DNVXDZrkfBrrYRU4XTtR1ALBO5WrDuS0k81U+5yls8ZW
w9JcTpedJOTkaItszXXco1elK3rx7WGc/7+wiCP0B6lvAX+Ps5f3bV6aqV2BT4crd/alOjgs4OHr
CobKnnAuj0jmEwgzE+r12tEZHDQogUVUtzblFeaizzsaMZr32KnpHf3KC1P6IAGQEYa1NBtELCrD
M2HkrYKTO/HZTLMxqp925rKp0JwkCUZLa+YYO2c1gh1AfsE6QUN8uj3/pLyUcQcLIOAv4PB6V+VT
9YAILTurnB+lMLAnKe9R+pyR3WAFEJiuCZJNLk0GFKLX64SGIH27ynfmfsGYZWRnTcObpU6lB4SG
6YAaGMqlfgURxExuUrwYS888VNQmI7v2Rf8aaxTX+hRK4rLXR1NS1PG6sByDcO8ZMUUXzNDP0Eug
TLtodi+m5lzahR5Nb8gBx5cKBNqo4VG02Ao8sE4lod4nNXrgBufhHvMDQimhCdnONRz40h1Xj1xN
IsUHpSxxLc4+eMW33VcW8/M6PUgY51J48Kh5W9iQukKfR0vmCna05Y8i/U3Ne7Wq7ygKCzUHX3sN
9nZzV28zj0SP7c5pG+QfpEyDmDLUjAj6bE6LgW9JWYJzT1ngO+4jcsvU9KzeVLahRIi99J0SG1T9
v2IXCd5ZjdC+1YIniSX21w06rKJLcAlqjQzMPHH5e1cL/whKw9j9OwblEAgatbMWz1szA8tFFpIZ
s2YkZGSFzji4bWCTKMZojEt1X9SVp4ObvEjigKTQLxQp21fbXbUXhVi4K/QDUvuOt+gIt5km+kDM
H1KJpzD8DVeAeCQbxS2X08HdjWt3L9p5aWx0jkGFfmy5jAE5dEztTYpGQM9aOsxAsTcQOGgWLjTu
gLVfGiYxwxqRhZzf4FOFtxOXzkJB7gbO8Bbi1TfqVEgVKJk1HrX1BmKTfTE9NIvCIk/I/PuqXWcg
BPNj/UrG+4JNAIHOJvBe+4IQhqSqQQ+x1a0eWGtIdM5184SC+6Rw8/X4+Mr518NkxpumoqFo0F3L
3hi7sZtANpvJ8L8Vzdf/3vGm1zFNnpGApUhu2SU6lP5ECGMlREfXnJyywuQFEjfPWWnQN/Ui7q4I
OSsPXP1nY/9oGL8eBB3VMmik3Lxn+nNct4N5aIsqPf/4v6bMz+039X6BV3UTObV3shXEhbsgQ4v8
ZUmMzu4euza7fwkoUX5pci1zrugVIwK2m5TqUOLqdtxiPOUKfIEELZMGr4IHVOAWNQ8/IZLrryaD
LTrXWp3GA0HucXeMbKSPxDijl+snHsG4BSIcqIrgAh94C/dStbh8+IZ/DBb2rYpgOJ8wZi+gYdYE
/rMXGR8Lr7/gpCHyrcblDKHhKQmvzvDmlpBJj2HZD36AfvNRKRFW4rITh/foEim4faTR07QPK6jr
cpX1cvLcOclYYIjXGmNgU73Js7lPxf3YgG8bXrpdPRn7LWKSSj3IOKwJ6q5kq7HFQVnrDitabuNQ
TToMUpVc12KsT68WumXkv93uQQ3BmkKUb4NoPnzBX1+6tujnwTJBWAoP4z/UvJjKdglisHKwGLar
GSWLM8ucHgMVYtSmWJQpPSQudsf8HdtlhrhazlHcrtpB1rzYysBgXN9ilQpKsL9HeYLP5l1E6l8j
jCfr82B2/zGADRR9GLfOHatx3h7DUrj1FRyCjyKrSyEhJjTvTiy5kv8eQP/lgjBCgSFumsEcTzRk
LryeRRmc75mHCnPwGPjOuf3blzBHUf/VkMmpOTXU8HqWZPOhH8VCHIfvIW+dQKvF8qFyzUXEUhWk
YxF0NarJhyNCh0KNIDA789yrdDD8CrZ0CU3UCPyJ3s77eYce3ZH1AjqHeQJZdWro5YmFJC6RwtPe
4jBx9i9p1fTXIhKFZcRKpoBEGzxiFdyX49HkwYkiXkZaFsMFpLegGyuID3olYqlOgMAM+JIMscOV
jUxSwJKr4lxiv6IMVTWengCdeI1mdxVVPShPtc827mUAuD+YbbC3lmIT+Bc5lUK2/mu2UmW0mejk
MVVPSg1iwGtQLFHyATjqNqaRXmyJXTV6yn8Mvhsbd1xp83mH8TcceQsGdyzmDDWqoE8pc+yIwkps
ftKAQt6GSwaDhSgZPnvpfQf4yCBjFx9p+RJTFnTWVmnSCgFUozSj5BYo61AwizgaBmXYIRa41h9/
e5jKm60DFWJblamkjYVYkJCeQkpT5yKOyR21P0TapL+gUK14ovit5xe7/4hoBEsd7Ta3Mf3lxDRo
J5YpB7zBFmylUrxQe8g852RQfQFRoGksFJ3gruC0vYHddQg/AuQOj36XZFqHyUAYYvvFUlbwBt4b
CPBIFFSUO/WFZeIINSFXU2+qz8ev/cmDm94l5xwRhgaCXPniMFiUrJrTwsRPrXRpalqe+mS4Vb4m
K2PKIevGeo0cJ4zoTB1PCJ7TswxO1ZNJXc6+81iniMy+GTXeDDeEbOwkEKh3p/2KFoUMucF7IE1u
eYB1g/a9Z7H/jfgdFvNOd0LI1YTFP0+hHNeyvUVJlx695RjpukbWYeGS8pYMzU3pXbfNHXlxwxH5
yqyy6gHTqLEFaPF853iPMSDphzWMCXqjxtR5frnPgKS6VlpucXpnkPJNiG1H6SyoKTiEYwwyRhje
AVteu2j2dOYjQqwQL9CAYwcyVrUnrZYxSKaa2UTdTmPsZo/j0nzwKbZsaILG3zgQyO55kDWgLT2B
d0pbdOrdcfE+nUNLLZDNlo4fkdD/K7OfDzxvC3LJLlkx3P/O3CdCwCCHK5/NoSeiubw/I2juHONh
8GG4UeKHaWuuU6bsumYh2DKyfUcBp3J9If7NAWeK5l95X0PcxfsqGBmIFQQk5suQBnLN8StqeMV1
7BnJHGjetCbKIRqb1BP4YHnREnU2BWsyBkO5pYDGlXqqmtb1K+Jcw3fa0hWTNcQpHSGLj0HnOBnw
ZZu0fzQK56tS3Ya5/hX0fs6OaxO0jk32NoXMUePpjhKVjRmNBNqmj83ikBel+j0iqB3sY8ZPOG7f
j/500rNfImx7rp3sQdUBIbX+P9KjYigNHsr9Iam3LdAhENVn4Tf88y8o2VRwODLiLRsGkcU53jrm
XN7Nv2w8Knr8b2vrptkoALr0cqoApr1Z56hGWLmeyr2+hzH//WJhHxxzImm3T74OaFNDa+T9H+2w
FQfzOFa8LJWVNyxuLf+yMP2zXCDfgCQc+JajvbqHLFhdeUb3OqboH2ZApMfeAHMJu/r4eF9PtRZP
ofepTBw4DrQZWboc2JQM/D3XcocCnQNG13JvIhNr39cNhS1gAXy/iLYUXEzFaOfAjXPIfatO25Wu
3OVWqTAVo2iY2h9Sz3BUWmplpnwBA7H5sZp8jOUZUURChsdxSFKQQDyzMbD2tGLwDtIkLlIUbuZX
mqt0bWy2/u7Syl3f68+tSpTQmTeAUKw1W5DVFxOJEzuS4JKwq4btaLdBv/KQbtUi6Bxi4hbphWRV
AJt9b//O9d1nVZY6VeXFoyM/D8tlzj03Gpz1Fu16UfVp6XZ44F0U9JZyPLxvp1SygqqvlG4ppUEp
BBahdI51y5QJNIuAlVen7+A3sui0KimXZQ8QL7GghbAEzajAd1L5dfZJxJE0tcPjPmKMDgd64AVH
fPmMUh5zg/Zldjl9OTsQWIbEJ55/gkCQ/04xm3ZbaE/0BUZqMh6L7TrzzHjcnC3+SWm0fYLA5IMD
zX/g6A6p9fd4FIDeHdLvuJTW3vOhEgzetGk42hK5PDvO9kvfueFrrV0Ei2DoORbrzjq31yQZBaVh
RsBFHd2WDyPbu3aWMA0SGnq36k1TzMn/t2FPpC35eItZ7G9dJ+bn/ozJ49GCFCIWFyckx9CobRE+
SmZj0vxEXe/yErOSBM2g1LFt+AF1eQpAg/IvZqHQFG9cU3xIr6SEWtfpB72b9x8g0ejizo/gkNFU
LElZB3NhT8A16to0juMz1MWAGITFqQ1rcvmFMd276lJ8zcTjCTO80rnRYwwBjIa4NlJaqciS6NTJ
38QCaUzF1A03/0gugggcGNk94k8Xfgrbrz1JUP3EAtj0V/CiX5M54zx4LWb8apIVf3UbVupfZ/qd
hyjqXgdSmmG2KhBjikeMtFqjqKVfNTu4b9wnUHNyG4IAO9GQPZYHANskl/fH9MH/WGVZjKXkiTw1
BKAHsd6B9uZF26GWLMmUjWvJBZbnlga2VRMecFXUJyKV+NgZu82qAY3PsLz7UhRJow/8Yk6kiZi6
gh+098duAZugoEjyDsaHVFXnWv60QpCgyPMxJYPUBtPLutivLeSqumYd1hQ9omKJ0gK6xlnlfbFK
DNuV+dzEG8eZzq+LF/W3VtJJWQFpyfR5mCRPrz6w0Vx0b5yuEUP4Yr9cCtcC9ohM+kStE1NZ7rum
dCOoroLhn73D/e+29q2WCuZzsd8dzQO4pxqq5+ylgOGf6Xq6qE79pCcZMIseQR2/lNUJMBSWMFDr
vfbljqbtkFQloEQh2QTWrZrHsrVtVJA26GN71wIbjOP99XFuay+QDu+qPDbn22QoU4QdWqOnmRip
KsPl4ZWRf/WVcd4rpwc2Cw8VKOeLN597W75RRhODDDUjglh8m+iGvKTaJe1p7Kwm2uz5CwJ8/Eck
bpdjhzEkhtHB5b4kk6BqZNNyFOBLmSL8K8fDxpFnWw5f+eQomN+wKo2kpTMLZJ5Sc+9z8pGP6eEi
yIMQF6AFMhnNAWW8L2GrLLlNF+cAj4owfitLC02poNXeFhOZcpTb9zBAfZtWN1pw3HPAr5lBX0D+
SW+CHJMnjiWsVkh6aQeYfY+4r/vH+lZs4mAKXPWMWZ322AcnBWykhR1REw1BK5jGbFSSUWV92XzL
Iszaza+N1qnKQHMAWQtsbXGPEZwpBAY7bJpWEMmwufjSGZS9UPJ4Q5+gQbR3gzgOdDigstfe+YqA
PkYEUSekSiPq6M1KjvmFTUgJccO1Y6mAsPI5FDQMmmubmzuxdc0gTw325cSsbmwPgpOvAx9xh4pY
cp9Ti5s6TKqpnmnlvx+pjwjVGelkf8yftw/SDQeLIySfIGk5AqET1G4my+kC8VCyDhKjaq3XBHvv
XnRNmbOPbnnWTVgB/45Kvheja4PCR/ASyKScuJiTLV2a56uZP3D9tsn0t0TRHhfChIufHfbcWQnv
ZHhguBGJLDpz1CVimn9qeyjvFJh04CltYcltIp+KRo6haXqUEFg/3lgDttaLvk+6YJCmcEtlGh0W
0NfAebtBAjtpA+tteikBNyFx3t3E+Nw2Yjp3DHlYPQ7laPczXJdWvkM/OmKluC401rnuC+QsdTUx
NJ6QvBmii3zy8/pl4fOD80SQHdLcvBYQ3F+fqHfmL1LMTSYCOteDRaABZOcelCHsdPahkF2IR0fm
W0Lp71yY8HUlSNoAHX4CZegOZhMpGp8PZ2Jia+V29Y0lWAj/7mCff8I7nyvFlDLadTdegTYoW1E3
5keo22ee9UlcFa5dyWI6o/vd/IKkZIYIxFcQjvWlUTJGarYEq64owxddZvNvj71ooqWyhwwVcq6C
Mje9iWvyvCr2DnZbtVNwg0O460K2nMFs9b9E7ZfxH9tMtcQOkdl34GEZhU70+iT4mZKD3TaLeLYx
WVPlpgSTk+dd181/yhHD4lQ/OaC+TY3wlU6iS5DjZbO+7spq9pDMdJWol6NigFAQRR5g9mDO/KsQ
SJxh+phXdUXiyRuY2yuCXMkx1GkPrzft5d6CMeGXHKEmZ6NeCuP3yyMyCWUs82x4dyMFxeYBMwdi
yj8fYzINkHnaJ/ofblSWvK6EVfq0LAqcBsQDlM22MCrK9R+MreiyHU5ctHDDyEER98XZHfacQKCd
pXNn+TaNEImDLW4WH9i+sJqs+eIHAZGcAY+ZPM21TxVIVarh3BoWVqn5l3ILS3LHowU08PfFFfzZ
x77FjYEse4UHM5MFYYhyv3hY9t6ISmZzf89LqcCC0k3mFhsEhfX9BjqfsqCR34BV8wIbUut53dyF
CFtT9fnx8wlhq/YXiUXCeBDwL438Cx8oJJD9bWuspdeMc7PHdwmkpVJWZs0nuchv06ji3rwBzu4F
3FkdRO3twX3XP00h8o1ZG485dH1kth0shyEFzvqRtU7b244RhrvZQg091xsIpyw30eEyoaPYJWPE
LeTspmCczODIOasU4T+92N1/DJOjJm6bwI8b8eWuzlxTSOaoMNL0gl2vjCuOXg8BphN5TRI4K/1T
YgxEsCu4D+mVNirm9RPHgPddq/3fLAOw+gBuW9UjSndYCY7ux9bHw654qhiwO45Nce6+03PwGkpm
ucj4feKO+SPDxFKjd1w9hJXVcgFADf30JMgqN9VL5wg2wx7D2+KXEUr1HZpVGc7KPbiFzjlJizjM
egpwlhvMeks6/vCAYdZTPIX5IqyWcwPv7rZEDd/hkdxLVmi131I1wG+HDPPgFNQOM5KjOUk05TN6
cEEeFmqWzKEvaJlTEw7RSIIpPOx9JGw4PkEYkBeCqRjXlRM8Gi4ig2VeTIEA3ZpnQyHKWN5nkmkZ
IOb43UPQJTsPkZ5TGxYR5Ndj4q0eYG7yse4wCYzoaga0Oh7OvT4p/XvL/Vv50I0jfZ7g5q4YROkj
ejW1olpNepVSEmbA+wLuXsjGIGETe3xAsAMTkH9yebfLLiRW83C1sTGVu7FIYsgmQzDj5QGHl5st
dT3nBfIkawjWsG7MwghQGgLa4WPQbFAl4qxInSxOEcSHPobGxKgfSGQmWQH+AaX92qgciRnWbBea
0frQxHIuzZz2a8IIKQG/9Gjl6D7ut4Bm15QId5T3RMmQMcYVZlwGXBa9KWkSkr5mLP9g8aiHY4Rs
GWxsMFJfYhnC7THjy9p1yXx7sAAQI8/WNpCQ8vTJDfAFzpnFQ9rRivV3nwlSGjrCD8hdNe3sJzX1
ACcQAnsssGCXLDcOMmgTtySMdgMo1mL/deujF898EDT/e1ACiFb1aaziCMA01GkGd1GnScOtMZZP
2B5mP0JCFJjRDD3yBJmGmaJYwZRr2NPBCjT+h/txSRu6HqUNLz6pqQUbsMhJ9SpvzHXqxOxT/iZR
tpU4NUCZifes1HuI02Xg+yR1+9pqjW+kBxfT20vIC8X+z63tkVFAyXIa92VjxzYFoGRnhircjTKU
4Zc+OaKDbLCz7eJ8Yhogfc9m9GdbPggrTx+IUJKjRW6xbZvLg2vTCoXD6uoBMiDjftEuOFOV9cYb
boKVhbPAIDVy79R1R28jFWN+++LJsktU8itOJ24h0NPm5TDRHVZLv/4eYcv8qnH93HxzNi9k8kAL
SmSRx7V1Nb8VZ2JNdq+LDjQ+ucSODI2U59F+2DjjjvHJAI8n9Ubb9Ym2y/r3cX+dBDsSwUdqUQlO
JbdzygDFJOl7RC/aHfYhJL2rEygNEAOSEBe9jnrDPm7JxkY4qR73k/SvrjTNQuqGdaiH4KRT8al5
1zBRbgA+WSDG/2+ry45hIlOif4/XcxcbeAvLu2ekW8uCBCJguab1BasHdWNzFL0MNJ6GHJwwkKGE
wdQQ1OmFpoEt6ZzVHfnY7RgmW1cr/GzuNV8nDFtIe6neShDy9k8MTWy9nXBJgYaVD6B0LmV+1pAi
0GFV6pbc8erWI6jCoKQxQJfylLD9CIvukvBJ3NSEZm3BqYq7xNXZl+PBag9n2xZhjWF61133+h8f
B+Rn/ZDpcG2SI2+t8XlQYjrExetcpq44uo/ufaYd3snsQlTnXzYQmIMxHT3MEBH+9H+fWGeNqmPE
5xG/jXeS30gTgaWM/JKFEQLSz4G9f8kFe8+gjEDu+gDmLuYHBMG+0rb3Qh1y9bvogsMZ6fMPGPfp
tWti6+foo23HGMmAYj8HsN6Ev0bhTFgWDIMnUQJx79YvF6QKmbsACf2cFMjmqrhnM9G7hE/QMs27
HmAADUcUjcM4YZStrdshtZ3W1sQmKf9iW0rBAByMrVIBg2wIRXW60Z0W1ksyfndcD0GyV1l5lkP0
C9nl0PPmB85TIaQXNCiDpQxPUzzGSK6LML3XHoXeEXDJiBzumzKGkN8KD4YWoClm7kv9QO8D9ONN
OtvstwEp3psLq/9AjTwb07lYQp+QF4+V/c4iGamxOP4c/DdOviRoC6eQz9Un6iqk3qDbG5Uq9lxp
7RqaaL+7+TNrHiwKQfstoF27dmhgxco9C9NPUjQm7pvaBA7eXepqdZNZIu0WFUHNRhuqFdgfeLdB
wsCT3LMkVx9O7tzZ56SyjZdG5sYrn88vBVhG4afxvZu33ogcCS2sWeftFWq3Zz8KYApsdftE7u6k
Z264sM0K9tM8l4SnlTbKLp8nd5wlg13lDY4LQeiwNWhFUOw3OMgOSCsjGGsChiF7rv4slWvvejcz
KxFo9guSuUpBg1cQIDhApXAjmx2Fa0zHW5oG7qdkHJa+GdrdpYLGQwTGolG/pvfROm9hlQIBI0XW
pUdmG2oBxS6imNgoTrTVIdRbo62XLKTk2HAc1XMSRdCNs9xFtCYr2NyFFu4qLmqF/8T9io4SumFt
pkyvxKoIFIgNNbQJJlXAteGCkpebuC7iC8L5MR9SgrDf701i8aiKUVeqHVVeOIvp+gGeRBiQh1G1
kDUVeV+yS79SFWZERkjyvCRRUO/QYa3J97ijCex9aU9yA8moF/Ypq4gbwRzs5Z773GYxmldDOOK8
eSKVMuNjT1s2BxNaUPm5xg4vZOLfzCMcxbMRPpbfhWMxVFUbr+cEkcZpdNZ/7j/OujX86mp9a5Tw
6BT1SRdW3T4dT86qZ9094PWMpoYsBWNo7Ps0QgWsABcucic3fi70zOeQf0r1ZoMrzsrAr5y03IWt
uy349RJhs91cJkMDNC5JdYy9l1pXovgwaApiivWmIjUap203OnMib4B9xlxJZj2XL/Zc+t4bLwEx
EVRACpk6sK0ENZr1Tku4fzS3Tl+7jwZNddTF3J/Wv8qLKaf43/jgdrUwXT1ezIi1yMynJ3MHkrWD
KWRPTKsdGRB3+/44GTTPGIHGSUL4ydaGF+Ye/aeMKzQBXDfvkbLqXUutHWwAse2OwbHvjM9bo+z+
sO0Dmrbx8cP/SgvDsruhO/vE/HA0dJN+jT8GJWf9x/RxUSEj1MuCbc+T2PpQ7iSJxt4WEPJG24Cq
0CNIywQG7LvvtnsU2CGVo/bogzAxxJdHTHQshNL0jnoD+c//Vjatd3poHZnfuE1cNVGDCcCKQY67
h708RmVxQdKEExCqlfnR9OamKgC4QvztD6qMay1i/qJuVm1bI3UExWSeoHio9G8TrvgfFoa9hSpF
ragsH3rKnirZTu7xVvajFQq+KceYiAfDeQBpcNV15aLYuoL56uxVQi4lrcOA9s2MyzK60HdQm3x9
ugV+bnBS3w6uh/O5LTk0xi+XtVH1fFNOWadeDHO6G1YoPjneapVSzZuectWY/kGgJQmnyZmnJCEy
YSFuh84NkJdlzUXBjw6mUGAjYyydM2VcirqX5bZTPFWiBE9xLrxOlgIhlnBb3JCVu6lYxnxhnkaV
mpCgEcdXQvtebH61X3DGZsWDcy7KvkGDvIuH5NblQC3Nh8d5uynyA39NvI/wuHRpw2QBe86czqpr
WPBnEf6qNAyw0M+XDGUdNFfHJYpeAhGxDcpmPnNiJAfoY6UnVQtuBwY+p7bDsrwUmeSDsgiKVbOU
CybixUM51o5FQPMdWKtOieGuQ88P8b0eiqLQijd7rieOY8iii0ZAiFsIOO9UN+Mx/bx+0J/Ick2b
VHZZDnq7QtwzcZslhEQuc0h2GTAZFlvf5ACe+f5+bBinV2wzolMY78DbHPeqh1mxuZUwShLyRPsP
h55qyUYHj3pQd/NTS65MCAyCPOPCYOdQBMiNWNarVrxxavYEYDNL4tqpEbi4CD7AxAdmNODHq+3q
PUooQq/a1HPcyUwI0d/XTuaV89DhT2gn4fvwGYZnP0q04M9u/yQ9HgkYpOSta223Z/Ib5LGzau4S
d2EHT01HfzkAIZes5ymZBMeJ3jwsDflJs4l9mpOpiO9Y+VOMSAXHcxJTVReoZmNQgS3+PMU9WAUs
ufgYGuhi084VNyERJh3MihO94rRaXpXi7UlhpgMZtRmUW/+aydfywfrJ/hDG2hSqWvMy704lL+VN
z6qtMQgWUANM0Tn8YlueBmN3A0HrEMmGlaGEcLLWvtJ+Mdpy5s50VwiN+yEh7dBKwCz2OJ7SWrxn
reaxgRF5OEEI4/a0SNtdTDzGbPMCTrC/J78RsKuKUdJ9yxU5SKBKUMxVUDQWCLYU3yqjX3lzNvOw
fuppRNDna5Sj8sn/XCLb+N+7K4rRu9rl25fQZTIhYTRxZx/vm0BBbVYy12eHx8Y++DIdE/P7ZFWA
hr9ZPPaMkEdoYizS36pzXD32mFoY/lS59xCH6+pz1TcTc1d6hp5vkNT1d2eIhrd6oB0bVEZvcJpy
cIKmqOeoge/F7I6y91rY//xzT0UBU1UbiQdblHhPzRNmpEDJse/MD9WA+y8RlaA18qfh53O+udHI
OUDOqg0RXRPy0IUawRaZlpKXJuds5qqYtzXNapSZeUR2jBjw6SNyXos9mtAWviJ4Q/z4UKoDvDbh
alEuNklJ85a/PoyZq1oEppWz4uR0R6h4lM5jMLV09m9asW/WXgpkl6Kar3OPGrOvHzp/7BhvvwDG
71GfU10OvbrBo431md1Lthi7MUbY8CML9CZLbz0tElIi57jPHkfYlRMV6lpLjkpo5buVeMJS+zqq
ZaLkE39txtniyhLP9b6porjg8ao3NiJQXKu4gdWAHP2AwouYVUJnbe59gXt9ly9hXjIhXkJYwfmS
H7FBCnFUdLjikXonMjb23gBp6z2IqIehVA9BxhAn696JvIFHOtaV+QiyU+kvzsQFQTn4dtKwTAue
g0pqKrjVEl8ljLibuSNdYMtYn6NHtOdREolYAsyCQRAhegWftcW+L7uCH5I7+UvZJJ+ztyd9cSqn
1QIUV9wv4BIsdeogspk7nKCwV99cySaJeOpL1nd5+iVGen59ZkQlUTu8QywLUbtk0smZYEHFXe8X
ABV9YcQXyknvjQxnVYGuiAOb1rM1Dilbqx98UvP1QpwHo6DxHQdzyy/a8471XVHMmYGEnPIkYfXT
dokwlqFk8+AYMZrg5SSINzoruw9xNBodQgVV2OoTq4i5pNjC+CeayTYV0yJW1FjqWKz3XmY8t7VU
/UmxVz0pqrIjBowCiYnRyyD59QGGuO5KwLvm6pblSGSIsPUdU1lqNf9q1e6l2BEAK99AGPeNr/oF
GFZCNg/hOsv3ywiiWNMiuYRXfcGkjPA9qySVjIM7v+iQUPXfDCsjDH1PPLTa1Bd6VaUG/r09VSxr
2eGis4EGAmi3eIS6+iqieM84Udx3ZPbB7EBJfc7sG2dPz56pWe+5MHnbi3Zv28Yx+Q4lVhZHJ0D3
jzch5VNCBe1TLmeXVZkFw3xNX+hqnxV5EHgSbZk9w6z2Ppv+vBI9wtHdn5aAxnIl2TOh7L+aA+2a
aPVn62imutNFt0HuGWPkWyd/VNEFEmBa5rqL6mD4DuNE6gooPEANtKxBoHfx1zLMsHNvr/YPxM6i
cUoapMFCYn960PRFCJYJ4OAvXkArUspywmPh7V1lS8fHRimsubOPuyI4DHRyMFGHxSddNoD/AWxQ
y2OTINjMQqBmr6N0iYXFkjj/PO9kDPiaqDp5yyAilTbVG/XrmDIBDRG9FvOgmxMT9VmNhKM5NRQg
hNT0kYnmuDZsun1e07STwmZjqz7WH8O+u4nRKFvY76pcBCEkw4RFfP3fqeft+hWmiUs0JXQdSMo4
Vzc1x/HErQ0FPlJOzdkkmwJS6TBz2ob/O228c69Vrywc2opy4oFC/qI1SHZVfmsW2NRkZ2nehpG6
eFfkP0Basn4rp2eHv/yHPAJyYCSVhsE9XxWUdsly1kYyDioK5ryIgjbXHpttqS+qa/eu2ArAJy6r
lvilaWEM2esUuajflhc/BWPel2RH+8fostyyKJGeZxrDL/6GpVkoquFCuIy6zTGw0R61nwMzcPHK
ga3m2U/zOgvpCKnvmxqUWeanunsS/3bogZNVQI166S4Zj5SI4fjCBkoBcqgz+I5Z1WojiB+dWoek
YPbts33T4hpwXk8X8oOufToF3UYz3z4L0hPjW60QFkXQnu0Gh6+k0se3leNm3Jaq8K0P/HtRrhYW
qMhdVYZqZfUPQuyx3KDoA06WvrnA5RFBZIN+B4rug2sKGpk/Mk/QCVHTBiO4gz7T2XQGgPkjBc6Y
pNnlECyEoSmGOiHSbKkMEjvihBa7Csz6f8lZik1FC8GvrINdX9gQh2fNHX3hw//u+jUveg3v+gGh
vZz/89w8Qj4FJN1+0UEOvAn1nkXjx7KeVG4GRskBvdcmLKUxtR/gsvTOAF6K5hIQ8WPS7HjsObv1
xxAivXZKBmMOwrkDJOuFWE2faQWyoK3ncbsxgGut8EsmTJAgap8PJCrUbeRzyqLQIb0xMYTAshjD
qMUyURYjJPurB3RqcuVWvYdoLkOuMI2okewAuPP4947RnBUwszs+ClREO09k0REO37f+SsuyBKvg
8dbhK1JD7hd0nHi4Oog7jZjnqbupTfjNjVCHT5Iu7FxAZQvFC8sFuxH4wtdkX71NXFuISS3qC+fy
SvdF/K/aPp7P9lcA7mh0rqkXiuovbMvyDCc2yzlmFXNyIlWTUgQl49ISgrV8I35Y8UeukkQfXHyZ
Q5YIQiQoAjcO6RGFN7z1zLKCbRcNZ5WvMSeW3cNqJO+xG0oLlN6SYF9/Hwis24U16OavFKrO0Fjb
Uw9H/yN9YTchk/U2tAjwfWYCi3nCWDFyiZhZrFhD6K4sHKTkfYN6txx++aYdiLEc3V22PJhB5Nt3
rEG5qScKn6odrby0rL0nwDAg7i+fWIdcndmlGwIDCEm9WRbj4X0+FxIcL47C1fA8TMYX/OtxlU/a
zgDVcwBjmHxMdkaxjuHri+9UmpuPBOrLdqg+m7zRs3KQ5UkI7V6/epEsp5pFQ0kaQxOWrxQJS3wF
cFdLyNPwXH4YNdMMzIGhnGKmbGI3ja3S4/809Dc/I/UUS2NqetvC9Mp+RhHfsiSW28zyaDgP7Wny
+QlscELEE9KraIUcSNx0F8V29JLd7hQ45e5LeW6tXGeSral1wvheukPO724E3F+wByVm+2yF0mk4
7xoWcnUpVWp/7Iu++D9rGvEj5pA3rwP5/tQqA6O1BCXF9us9O5r4VVosISlDiZG30dGGjN1s7LoA
JsqBUUtJeB1taLS/gIcewKmr5WcV1rcIHhIHVdUlzO2H+uI0y1urDuIx2qZRkNa8Ssf9UZVxxXUh
WOfNP8109JkJuVqVKNQIhGI4JTMY8ZOnIBCMSyRyhx34XTQQ1puNFZCfcL49OCvYNGtHZrqfBKVP
pDLeB+s1COhbeOGT2uEpeSbHzxmqL5eo9hCKICpokIcjrBwvQc97F8uxzBVZw/qX+qwuegjuRzO6
NtEUMKFWmzbG5tXv9dWCy3p5Vl/uLoGfeLwqtdFd7VCfIU+eyPSe0sUUGtbSPF0m+8MQdmMbOizQ
SYBbAAglxIPdCqNtE2M6zcifywzZpg1M8GReNBQPj83S/zAOM+Dnh8zoyfeObmBrRNTQ6/8iLtYX
FmjZ1yQe4LJRyofMUKV+aoGnT61aVQuVTI+nP4NJJBcmsAjHxALg1VvEYtfyhFz/AbuNSgWngjv3
tnCOZU9JcjFXWUJkLcLa2frOimJpCEKprP36UPmnT5etz5CRgR3T0EQtyS6u218k8oeUrJWfyg6k
sxdyBl6cq09Me7m6EuzDiOqIkcE4Dwd/ddehCohoQ+7g+DZZcxQ1JlWnOV7PJLife7NVvHuGl2fy
vOv+NHXAi+yfvYMxJkwPl5AuxvWsoFWOFAdjHL91oWWysToB9sQlzHR07hb2aUx+MhosKvfGJltC
hweGFf0gIGHlJhk0goWTKpLmxut526x7TowUDS7gXV5datvUsAkKTQu+KnHSY/9X7NHXfA/maKtS
8AuzE+r/NTbGMzE/Fvyk+qeWP06Y0kQ834yyCBSeRvgOJD5JQgCS61RSUFulaVaa4OZNelrwGb5X
+NArGEgnRWPDKnQdpwa4HzDeBCT7qpZxH9VcmcbKT7G29gUbO5ODlLYbhtFHofiV9gyhJZ9etziU
f4rqfOZVI/Nf44AxTJaBiEPZJ+opvjlEQv6ihOV67oP+Wp7tO+z06jLGRvo+EHhjeu3WRjidfyoD
aoxaXkPYwCOKTEK2yXDt6inqqWQYMvclJrS1GXQAeOaHfR/6R0m8xfXqFvKkcvYe4WQV8u+jY8L2
0BV1kecccdYlkIUD4HlHtMpKgxyrYqLBP66aStdjG8DTAaFMr1Bhko35+TrHtWdjcZgzOhIIdjWf
iGinniMcoOPEBETG7iMkGLs7GzYLLxRyRCcjOK4Px5nq6QP8veqbsKJYoK2WLf7juwkjFc1LC0xR
MrDaNBwkWsfJun57QNg1iMH8GCk90QDzykeX2n2cpwi6jJ9R2vJE/3SFdV4lsb2tZHCstvrp+iMd
7aKazFDJO0Sf8Fi8QyjQKHiKDKFvaDE1Ta3scJ9Es6wnO5c8f19w4QAHgDFb9uKFkNNOgTQgONWc
IurI6a8OP8/XpJ8lrhhPY0o6GAuSrK/U/OmgQbNhyb0YbdpraowAner/QE0qwbpyu3aGEpI+MBwI
CMtU9JcKnO8DmXnvLfKTESgO3S8njgLrpquugNy2biwAP8mf4IKjDowpYU4uZHgwWJzHdStwS66E
49NxSk1cZDRtbE6IffwhAC4YzlZSyV5Xmn72r2gtJVEypJ6lEDlyQ78x0nZYh3Y7E7trV+mMbFTu
7+xnV1mIdvpDljz4gCOy+G0S8rjmtOhOIj3maUJOML65XJmrJI+dSMjGw6oeshPVngBvEC3uLfcr
DON5LlWhGpKfzEOWQ+e8wq34VmkNzOE/OBom/KTgOCrExfrVyEZ34H56DKkR7N0HJqgKMK7qUmJZ
Foqkk7l7PnN//rH7BF+P41PHDZnOQipOuWGrQ4tvn1uVQbWPRw7dTZAw2P/EEpT16gPaW6//yoOh
o9Xaeyscw1Lv3K6+11I1h3c+YaWvbpaUckBjaT0lkDwrAwMN5h4iNbMG+8tBs3jc/zIo+0Z1hdal
+98JPz8GYatUp/lEtrbBB6mD5sx9kNc8pQuINVd4t1cbh8Tl90g6T2gO2JxIErBf3TbtVpWdvlyY
plmLHMs2JPMayJ42c+4Zl+GsQ5GA56Sj9ecybRvp42RW25FFa+rroo12Lp0cbX7s+xNFMzQeijGU
V7suCboFinGH3dRTQe0xXCAe+dkaFsfUlIbxrC4wgK/LUHL9uP5aiQ7DXlqmxyO6nA9qBSPqJLfc
Ilkpb/2qPRz6J5fBfX+GquStgONa4vsirYzYczRaY+VxUs7yvWmpbpJ6uzj3gp0hQtXTpqvzWzf4
uAEulezARHEkBLPoE4Ip19upjQbVMEc4xy98PNVfIIK3smDgDvWUnhpM9ub/rZ4o4ZlxgoMWoZkL
DUTvW4TBvJmBL+KlTM6WlVD6idJc4cl2/UZtd5j04TqvbNLmJ2eah0vSNbdrN7t/eDRdL8zVkd3g
uLr+nC2b4FRvmogHxv9gZpXlZGI+IiaWFXrIyrZlevMj/6wgHz31qgy3c2xsJyNCkYW5D/xi97YC
JLngva+DgvU/6ofDEpcyXVSuIlpkGUzTEXdgJzARulyxI+kLi0/Zk+FPNYhAHLrfNpHBZsSI1kRy
A058rO5qE9sZqPJJE69yqnAsi6JCOUsr8DgQWXun29EROP51q2HW7v5Ear9A71nVVEQG40GCFSE7
CUXxWBhNTM85P6nneTVe7GgDV/vzfvU27uO3NWoT/gMWWjRWoi3M5x1M0zT2wt0FDmvAIgQaXbKq
QlI5EVsWPkj/I7l4vIZxzgGG5qQYHbfsr404LOq6AEvrocSYENXfZaA3VoDikXlrX34/WhF2Ed9V
AyIqR1XOfRAbmblt6HIc7U7s6HZFVcbRs0VJ7T6Fp0AhmQuCTSngieuzXN4+kTyODPQ3ahNtrV0i
/dF7el1SGuC740D48Qp7b99vkW8uNe2Iu0QgHti9qK61Rxua3bp+NnaDvSVe11ml13oH4xnEiupU
MDddSvAX1pCddVb7L6DhPncXq+I97IB4AN3fIctQIxbJhFxDVTVUrj85WH0Lr2c5fuzWHv2VKBd9
PT7kQ8v5TRwVOolyyFzXgKW00MQqWv8IRwr+pHQwbr9sRdKj3P2A1VaqA/JiM0Vvi9FEUtnirBNH
NhZ0vja/L1s0jpzOp0HZdER1liQ/SsTaZ+z6Ko+jLsPYfoYlKGsU2rLWpM75B4Ovmfn8T7c3ZInP
QO+Ldv+899x+tOaKMWJVKy/7EWnzpLaPgvlAvTM66f9cNbD6YjSL5FAtjkqfFBv6g0sKjUqxNNRY
qTlCwoXuPpNF+Qve5i7aV9n58oQGvKCNZobNpszh/aMq9HKOJmyEMSjDplrHBZVxcGooLC7MhRtm
ZNeIVVStrj7LHEEN+tfRrdYNSm7/BI/lg+qJB+BB47/qqmpRkLlUlYBHRq89nBCfZ6aJTGn6SeP1
HvxqpERMoeVHK4qXNHJZtSB3vYX+dTVVAUVxX/uCAYQ6zEeRh6nNXDK/sBoNlgPntWDXeui103Og
mELy/dMjoI3IV9oA7CHY7xvtvJqsMoGfP8ADQb6lnqNjIY8s6M6B+01B40J8BkWa98i1saog838T
srJiMcFSUh9j/ZE6rE50DQHpRpiM+MT78nyHQNgZS16okkfnM48jNq23dHO+EXRwcaaW7jKAizJm
ghtQ2dPm0VbLsijPn1C4P56ig4lGrUktnyszPmAuBusfh1UD5dGQ8R7AzHLaoIdo48EH/Ohk9I7L
nEEtGklXVd8x0GwknLsVITd9p3pgRCz7w9FF9XtJq9vl2yah8XnS+tf15D/uJEKQc/RMhXYyt5Jd
c5HPrpELEjMjdkYJC5dDdTSAzVL49yWunCVlHQy9oEv45HHWiBfwa+nPj8ojNMElbwJ8Q9JP7FAM
KgeHL8+6h9OYbeLByAjrFMGfq/0V7JXd5giHtkXvgJxvIN7sMRGctDeHEvS0K+7gxBxd+p4uHv/o
7sBZtWFfl0v0fYNzNUUiPxTrH6ttz3qMgyYkcRtbpLGC3UrhLR2tbN+lsFeh8q/jdXt4Q+u/UpGB
AJfM6FrFe3pFF+7YMWLwhs6kVoN/BJsPfEAIYS7+R6Z7W8valkdT6aiOiBTdsFgbt5bBrvlgpF/Q
e/4gZo/LU3leNfAmkm5O2sRFS1OQsgaeEUJys+qS6VnIfZdFJzs2W13jNJXZUI6+RC5JNHgtMgjX
aW5ESaiE0lAg5BdpHFulcCcnIw1hlPW5fFLMK3g9QL7j06gxzf3w5wpNqY2RDMPVnnQY3A4bQnRI
hs1IwBKvliVizrS30VJZOyEENZqqPh36BAdmfrSs8Uu1HHQal6RxkA9G6bOBbY/7M+BtERuubohO
DREpAwKN6TimmVZcYhXb+px+ag/EA79U/SpXtedC41a87QCCA5kqjRjDT73t1yKySX4RYUp+MxHb
erZotaBjV4rHRcW5COj33tXISmFswbjzpd5dinTwmUdWTKoUboMwUfER9NbJmyMb4Nha49G23BGo
wdX82WRlWv1nnaAab6eAsDGZ79sEy3AS3m5rbFcSg90z2gW6/NVcjnFbFPeQVqixEdI1DjAigRNl
qobT2VSv18rJxl385jN85uoRWEI7u9F6rcn8W8rCSRQqe+zgYWZBOXDFo4r1KA6UUiQLl1ynSK3B
Q6j+/41msDz9UyQT9Dx11n7kh+ya2uwR3xpkM/uP0ukjKd+cp7PsFhK/Eq2y+iM2CwSCMNlAnUuf
tMKRwrmjNlALlLXwpH/95E5rDVb1kLtatM0Y6PqjaYNX89wZ43VzpufT8wQToVFV6tAWEsiDnINX
Ew3IRjXcq0au3Bm3mxTi81reu7SgV327u0eqJ/ZGzZUSx/DjjgQ2jTh//vgmevO6QDJOlbVifVAR
piZJGUdKf3MrKMAyvO/5ezeQtTezNuY29UnM1j+tA8bPnGfHjBjxb+/9Irxx1wB1ssQmZC2A4MqG
KeQIw2Tt4iz+w6+OQkSqZF64KFIkNbkm/l/2XhB63t4zQQ+Wp8MkU0G56koi/F2/7MSSedQIghZX
z/L7FRXF8fwrncHkaHMMjaCRDRlMov24HS/3Q2RMXfGhdLU01lLtyOaxClcV6smR0TOteZvrGMGq
u3quKUORjSPROfGb0Oaho9WoL1oDFBBR3XAxzYIHXVly9Yr7DXXhF1JgiVISuL795QifK590Qiq+
Iv9ZbDJAsfpvVPr6gKH2717UxeOYnPaaRkuSQmdyRnnmx+5USK5ZW1q0DRz3zQv24/WG70B8TMKB
bfxPujYNQW7om7h7PnxZHdq4rcCNm1htxlVkRIeOa00vaLWVBS1+OPOXYx//Gfn7xt8V3cyJSakp
j3qpcfTfVTK9lTpUDYTg4l1jVXcVomMYpZE2s7rpTuNtiH3ar5tVW8xg9/MZ7gl5kMi0k6ktOqu7
xFzqM4hkOBmoqafu0ab5PS3ONtMPJENDtqGmtwUrEewVqfgaGiJuPHFCWbEAFI00DG7cYtbo4LOO
C8mHxCpwOdYsj1H+2JrHeok5whAtgfB8RrPRNtAHUcmbXiW0kMQwVmEZRirqKyd8Dmr5ubxvw8aq
h2mlqSYvygcMbLv+L7M9TR9VJjGFaSSa51a1oDiAc7YbhkFJJZTS0fqSZfaLtaCZEiUfKjp9gv9D
mnGgckac6jqJX1edpsPHtlZYxkDywTz/k0elOtlqx3HfJ8d7RZ+e4PL8xce68mSqxhvcz5KG5DK7
9DJaYGoR257/PCfdlcKpAMsIyUHRdI5aGssim76jRlague23ytRL4zsMvHbrULp7HqnZKvjKlkp3
j5/HF4EDQTWf5MZA3Q9QchyIQFXhfHW2a9b+RcqqhCYstzflYohQEhGQRJfG2wre0PWilO+pAVWR
GQafvvQKkvwQCgiXrAIQkPe9J9kYWXb2U6VFiPq7Mi9B22CiI0vthfADiKwO9006z4r+qDcBAA8y
aQAzSp1MqBmOtADVm+GQpO/TXJDVuhxzVFlewrU1I/DlHHiAqA4UoGBhdYVV4m+Div8a4P74m6GQ
BkrOqauYGvT4DAQNRM4BsBooKfqoVmVwvR3R7pBUQ1GYCLT3HFxHOZaG4njaktE0v0SeyRE/pTX6
yevBzQZQnkSnqZNI8gnGcj64YKSkLy6qHX/2nsXXiVZvd2qWGYXUFt4WoVGiuDLyAim/Fn+LQ2ql
UPcvORZj8jJJYMAVUZqEQxDel4rPPtHovse2iu7v0puLOGFLpXp0Trvq6+4VbHUAfXVOYs6ydn/O
Z7UNmzduxjv2MOFNHtzjcMb6Ja0VaYfOPdujuGRC9xB2R8hnWyy1FE2P2XjDpD7QTarKcf+2Q3y3
z8sEQVFId89Xv6EIuZjrJRgAXpMlAO9jisma4R8AtqSSNA3RffVufhuyFCIqc9Os3jiOkNjjbb+S
u+KHzCs7zUvr1jHlkzJCarTfgtEO0e88l2j0yZgMqVNZS9Dj0WFyKchHxtbo3td3FxSj8jE0Vn1x
2pt3thJwxjbSg/SclmpA2lqCLkwxo20PFWXbz6W53sGSVlAQ9VYOtyJq0O78ei+jkH5pCMYddTTm
BiEEAzYDqfjwkTmNbGlmtwzbeBYHfFdKLcl3e7l2BDutWpaz5k79KAAVpOF2jw6nn8RnRpUQs0Rf
OzJ3cadtBFwf5WROziAJwm4v6WoQ0EQK2iyyE+JlsbeB1D9tOk00ZV4cRkDHNjOChJnX5+0qMsko
7dkzgvItw+ZOtA5tPV+QVboxYt+XY1t669zWGFn/4NvS5+JOCNK1iTfEvrBDSKC6E+PL5LHZhnmR
iOgF7Z/jPc7HOamI7dJdn24EC8vd/rp0sSp6l1ykLLQsaWV6Tyc3BUETMDL80rSRO4NMEiuGJuBH
K/0LNRO1upzXkCAhTqlWeJ+yn8bauSjCpQzqgA/CG97O2CIo0LAkeUxuk7mGsK0mwXLFZqFvVANd
03Ae+S1P6aYmhL1lXc3jq0neVBYXlVnF6lB10P+kMeF5+wLxEWKaC1+NPqlLDzfh1yCsu3xFPzYu
ieR3VcikFJnjISIDZXiRX54Ye52Ohdu1PDgWH3izfdpQlUutR+6Y7d9wpARKCSLhthwrGZD8I9a9
5YLzT6EZE0ZlXjtkXYYcuDpbzhB94hlp/R1v5Flj5Onxu/V60e+NXmrwTjAs3jtsqO7zkNSEj5KV
+v1Nvf3d9QBCFZ6tIpaCp3+JOqim8AJV9TEsAMX5JCBIVrxqT6G0b1N/uxMPbmYKp6Pz1YC8AWQ4
XLAtdigOJFSGoAfb/pwtAMG0zMXwyiApD/yyjHF9JyfkE6S75nfvrKVWUN1etOKUkvGQ/Gd9Q4Lr
nXEvHs7j/5CmvHZbFUBECMWPs5QdJ8tvDjN7cMOcIfigSrkLhFwT8x6vEGQEce/FX2iDDa+rXEvl
/Y8gdnZMBjvdwqe887ZnMnK++t3CvhTi+rCO26v5bGJCfwni14BQX12VeDiIz8749PfJpeYkM1zV
pDWu1EJ0Qd5+i6k7c/7MblvPAzU3t4NVUJ2XyDsjMzeRTbaGkiBStWZmBPmBzCpukFpzwTsFZU/q
ZCC8wf9DW//jOf8X0IG5VkXC+EQ5emrxWwdnbVcmiO81jAIQkDr9tkgXu5j6V40MKeuZydURI8pa
uhyn+/TY59tpWpHN355UOpMRk6yp2PROey667B8IoJeU7fTccd+2x+tIkDpICkDaGUoRumKNRYdW
sBTNPdOlISP2lbwgekeD/6w/+WlFCuaio9EjO10FDg02/ciV5uQi9LuSOfop1mj2KaVljavorWdj
RlnAv+XsWQrlzi3tcx3IhKOayftp684hdOIfkDZUPHvUBkKFWx6xup1VVH9c/16Zv2TNISeZTGXi
6FOdj7athpORJKU7NJwMkUjB/TIpUWjmORm7dmAOXVfAZ0bAMCBy5gNrSHa7QrvXmQsecTBOm1mT
8VQA1Fx6uRelOD8RsS0K49UxidNDI+e/KpGb0iaTW9LtJmXZEaAvWBR7vItAoKuTTm9zn2FiXEcY
rAp51iop3tPs/+zC1fGpPKlC0AmkpgKWWdHILDrOjxkJtuEfserSWs/NKYcvkmIddMtmzI/ZR4W+
Ik05+Xe4XAjyGfNy/sjYSno5GFo/8q/ziPFdW2e+uCmE6Kz1jOJ16Vpdk/FRDFGh1G4f3Iq8TBPp
un9ZXLo2FA4FWRn5Jralj8YkyWyUiBE5v7789hAacMk1k02qim+EkDxvTBGi/YACVo6hwDKcxL/Y
+bvPLnzeBx9bvoqDateS4t3Ql8eoayrRMjwv5gEghqzgDdCzKAduw/c8laYMxW7uufKpOscLlAdC
W6BwdynrLddhg3beBJEvG+CiAiIP4gTEuCXgOec0LLP4p2ArBovn+suOxyX2SAszSn7X1fYezMuq
b/REaKFS1NQL19vzXOf+Fn/++pEXZdHUZAH60/RZurL1uTW4n5xZ+j8aDqGa55SydUW945fmLbdf
ZwuRaXWUR4tYQRwgB+CXU98gFiCcGPkgQZmYVDLntFlzOl2X4vDYT1OwIZNCK85t5nMk8OVgBVN3
VIImCkDKNLhDc44YT6CGF3gmcZah1TnEX2TfmMHgYpXXUrm4ySBY6AICZkLHkpOLOo/4m8brvHf4
Rbc3uktxRvj7PmYpNzYJ1TKqokDnJ0efpE1RjKDJ9aAjO6+R4JFHeQGXa3G5ptS4nUyYNKQVacEh
15KGVyUhafXdaVuy3OQz6yWlLa2eZgdwsii9eZdtX2QZ/jVi1GsWbQSdJo9as48lp5PmX9IX/lZo
5r2gICmp7/qfDU4yrK7viCSvir/dFsL1f1ps9DuOwBxVl4Vtl2ugS/IoUttt5Mdc5L5hLqWd3zrf
VaK3X+w2163KtD3JbHLexeReix/ennNM/mySufalAcBqq+1HMVWCjMyNKVj4sBzWoPpjBw80WFIf
A8EXpUspHos2C8OATR95y7+bOhA8IOOBn2jYwrHZ71f+OcsTI9i7RdCPSuSdos0x6bWBFfofa+Kc
SCiU1zc4tkcm2gZeGvYy646tzEvdLeovoe1T86PFvRTgMVBz+tPgTmUpVlXTj86DCFIBOUVAIYqm
KT39PjvG47DSKFmolJpPPYFokw4UxaiPp7YSEkoJWJtXlFAmNrfdYmWTHTdhhKT+tyB5Oy1hTz2M
CNEU6McA/9Y6sQPHOW5bu0BuGY7BbPvGVFb3Stch3vkoGWbBhmkCU77JxGhbO58Nlup/dY44fz1o
umHgMOTBd+QejeJU+Olrhooy/W61Vf2hLScyhAybillXbwobOXrse/c/s1giWR/RI3U9ZGuQ8dQT
ldiYWVnsDFr4kyB/7R7QufXVZQ32ujrO2/U6M0Rj/wpDyqflsa9S1i7MezYktYuDvZNMie0QB7bF
7xZ+EVZR8IpI0q1NSxxLx+V/ZPrygT+uHQM8MlS1FkIeVv9RJOPJyzDsMI+ngnSgpFe5nycMCskF
RR3TOi3B1gbWU+20FXZ5/C7aSx8CewMEp+r15gIMs1DVJcGSi3skLyDKxcFOjJ7tHQG97cAP/+di
RXgmPG8We2/qR/Wpei0AMpFLRs8SEkqBwp4cZ1UmKYTUzrDEexzGr4DLic3x7s5acCyMzSRTP5UR
0Zw5FSr0oSmnYK2S5MjzlPwmRGuLmv4BBSOyENng4zvJJznCeKK/PIbLE7BOfWDGTvnAggDfGcsC
pEF8bTVOMVuJ46mddqpCOmVEGrEy49O2FdujuYgAfqbPujM6Vn8pI7PEakz9S4H2Qnwaf7Ch75MR
McQp/ayW78mqsPM17EMilP68Rv3kbpGPMFK+xDLAN1HH8dokAEEc6pwZ8H8GsTw4aeZTIE8w/baW
jjAnkQMznsQIbevynHcz2IjNiK1W0MYheAnLoZQa7u/5ZrANv2w8oCHNNbxixe42h4JRltrUm60l
xZnMjG4C7Jcbcb5AEOwIoxPL0dlnbS5Sf4fD9Bg43miCEWzdRj2qGUTpWjA4AhtjEI5rbGa6e06S
K+l/Lb1kL88EzE09Sl6KsNOJSLmUPrrIWCrPHpeYftIpzYKox64kg/Pv2/jcP2/Srye51WsD6fUL
N1CCsMMf2iD/MZrscVMGq7n5X6a/eDb3a0eDPOvSwqJ1q1JJHYwBLmkfwXn49DvP3IMbLOrQNrQo
TiNjullAfkJZWZ1RAwCqaBq9+5Yabjk1pVLVFQ/An5JpKsUQefTiPsY/4zauWfHN1tFSDxBbdVX9
xMaBsDl5OJR2ChlQxsPxdiP+c6Ur8haKBVe9eMX+BngJK1eQs4wmENHFBfeGWxC8808Gyh8gcONr
jyI/ZQ9+3nG9+7s04AjBEPY5uFXjrFuf9Edsgk7iLNU/XQTp2nnZG1UfR42FOF5nEHdQsyfOzlRU
n4hDoRCyWbImePFTXbDSCuExHQSzrVa0WtDqwrt7MbSg5wexiKbdHfS7afpwIR1QuMYZZH+lGVAi
aQOMNJa6DXola9Neu/fzlHwkVmCQK4hvLc7sFTiaW4aDED4jtTPkAKoFJqKvZDjpt366lwADaYTW
EsUtR+zLldW9gchWQpPixYOejHKQfUYIYa3l3v5TnUKGejkTTt2+w24dEfFmCvo1bPoUzdJkKmn4
z0gGu2Oe1rg40nLhZTwUg0Tz5xBbA46g4qlLPGY34kxyHEmAs2K546+PG95PU2YUOk0iILf4MUK4
uIJEKPMCbNLsOkuDCJsuKQgbuDVVK69b6HPZXEnQHClTnBcSrhcgUl1hO/QbeCSZPlABPBJCWnvT
5edmO7CnQj5+tipSiPEZMFQUf74c20EtpBppLdp+N/zApqhSa8vfH66sSDqCaqHRkfjZsyjjByuu
5fqn0SvDoJAgJUsw6aufrw3I+h1pmZ+5e+a8vvrh7yyMivYmsFQJeZkfxrp1X2ngiXodqieQ+IA4
2O4ENo8k/lFjbNcQR4oGTFP/+okXMP149dpmrZszOGeVW400+JR96WxPal7nqNePPkYIz1MsOTrb
piqHOnsDTxPgwlV4PvwzJAMtp4QSbO0T6KZrOTKOX0Hl7D7xS2kUfiDJSxnjuO+OcrcwamGkPLGb
kKvmacR74o9yr1yfQPa2pVmV0GIk+38M1l+Z18K9Y4bSisQbn9k96K122KfRo5KFK9W0fpNeU6g8
7ZiMj8ZOF0YE1bQtpBIJzv0WqAX/+5c8YXFwTX7JkMkibO+Nmvwy7MF/smd/e0ykVwFK4iFc46Xx
Y+AEJBQwISc2Y1xSZhSz9N3AWCv9e7DNCheC5KHdsjk859PcflW0gaIXkmoNh0xMbOcuGirzSRAq
+ia6AxtpQ2IWFspIwtXHt5asA3vMSLONcxQtkLfUEJsflsUL2S3KUGgBOP/BwmLd/J1vrL2vcj/3
avnt0Qx3GcukWK6YdntijLVHb0QZ8B5QlQ/618NPhcngUCmRPoZ9w8+Sz+4gcN0Uy9yHujZ6TQrx
VOCbF3v3j7ZAfJ9n1tbXCjfILTImI8YKcxtHhpBCny6ICicU9QUjr4uwdsD7LLg7HPTH5AYejZP2
WEstGFdyzFGDcYXdfAzu/Najq4wgWcA2Ta3JxP3bc7t9bEPKDIDqUwQ4k6mzMeiLfgPy7SgVIObR
lD1TiVvUvzEIzWqv5SS4+r70ZszRAqdtLxKNel7la/4H0DbxTlbpaGcegieFpVXD4mdKIm+g2bjX
bwvY7W3zWacOoOuonkNPb44NrADiad9vhg2rIuS+HrbHppLrz+T/ShUrhrm052jW02CBcA+TnzCC
RrCaQ2YdVfA0teOOgbh/s+fGQzwk97l8DBT9KY2JACbYufPi+M0fXjhie9G25hUD6SDSEHDBBYMq
C19/KnY2PbBt+ULU+StxxKJBUASSzUpsnJexeaENzS2gFMODwvKmWyrOxfT/JI5OTWIXmyK+/P+K
TopZX8Fr0W72yc98tTYzYRRGY7EEDX4Xk8XDNdPDA1pyeqPx8IzSXttAf18+bwwvy+aCR6QnVBXO
5/wmMzUWIwsabt7JLbrk9vMzo6HCGT5E0zwQA4kFZUgjHt9/GAkug2A13oHK5kHy6bTBxvuA1wTn
RrhFirRBOlFNzvLhyVcuKCqkIYQkA1RJrUSvczob4y1suLXTrYOH2y4mNvOCqw5CQJHTXZL0rWAu
vEPCKFs98PG4JF6n7cmI5tNub7bmOyv6hi5CmPFIiubur9/NPpdM7uEdXNEe4CMxw42pyPZr/IXe
uZTc8X28OgSVr+8Nbgvw5W8CiwOtQzWV6wOqZWkd+VTDdIMG6BO0nwt9UKZ9wDDh203gW6g0o1Nm
gOC9YZPnXwYGC9ynOr1RWGee0k/r64myEMOl2un7qyWzDPMRYn5CFi/6JtbbVvjtrrqhHbCIFDb7
rK/+QlRPHVKph/IOkA9H4JLRsEx+tOyKBD3yw8hxcBQusGpmeEsxt/CREsPFQ1M0QIFhxaWuYlI0
f1uEeQ6nc5wp7+VEnD1Y+oSuW7zyDk30EmVMdJRkyaBfUqt3As5wC4WWQbiMsFlxULPeGdQ5qet7
8s0f1tb7ClWl7eGyTySyrN7SY6rjluxOkqsqLc64GqIusG3GyEqX+IojvTv6gD2Rhw2P9sa1E1mz
HjdozzzO4Qy5cLxSUDnuYkn5IA0uBrPmsfZ/8pVulmk+Ch0+pr7CtEy7D0l4V0XD5ZL8iYX0Dwf+
DzOFmDt3hs37+kgr9bH1hDXzLeeKhHyPcXVLAEuzfiMsdNzzef7kUgvxJFIzT2znIfir7+cr06Bz
T/i70g0d+eZaUvu72UUeFAm9bVLTfq7/uxcZZKkEzs9CqQvr4Xk61QOJ9PkeBu05rQ5A1rZ6h2tR
bZtzVLwpz8uywN9pri8NILgllccCbXqK2T2QFzz6gM0oLQ/TTMum0OGHeVb2ECX99UUrBAcjE4Xc
i6TJxiDXfJgkCzwQjp8x0kbtyK99wyFj1HE6S/En7YaTO9isaSsV1jgkuH4A16OvEAjFsXooJHrz
MZr7gZltN/gMyHrvlSW0JuDeGOxY0idhKANaWPKkXwXvvq+2Do7u9rrCFLUgLLFiIOrP64Msz6vd
95usOU6ZsvnLYqNnLJE80jv+bLCCsX5NA/M+o2I8Fj1l/MBKSKeREEk3q1zcqplnIQpIpitcYni+
oupXQfrAD1bXk4eWUINY+7psxwBMHKVmCZDZv1QY9vxBLFrDfRqyYcZKqWOb6cKXgCQm+Dl3z5TH
1QoS0h+JXdtcEa2xfeMeygrf30wo8N2sKqycnT2s+lSseAnnwDF13p7j8SBG2wVvOVHgxfkVCrPO
CLH8Vrz+N6N316mXnduZfvD65j1xSyQX/3Qx+SwMoX3cxuToqT4AOBzqqtbL+qeGqyZ7muBjOnFn
BZGz3RPY1sw1yNwn+V/onfWm3Dl8rbcZbz7rm/UtAHimei1W6XfjuuzJlNTEzPSDPBVyAlMaufZh
8DO2CvbEkbrh2amGpcYXpJjAJfD/mMGEqvrDjwroHURnA94csEra+K4JcjDZJ/i+jOzWt+rR8Aid
q7WrsgX5P9QRp4VlY1BSTWhIQWEP8x0UQqZT5mWQrmqGdWmnSUkXiBtwX3cYhmc6wvYjdrCIBCHo
HeuXPN2HUvTMeWLSS3uspLp7FfAYkjiTwZZldsMRk+c6qHi7im+S1l40VMfHDM+ylVW48ujWraej
gZa1+OWzWLtDz5a9wge40s3XiEjKaDfuHsptVOP/lTinFlfIuUgDbgEOoJ0T28S6NkNyNzsitIm6
nltoRnfCxiSAjL77NALRzgEf/r16ozQgVrzGye6BjLKAlRdvH6f7JTlGR3Dm53D8+AgQGJ6wqWS5
mYFpKW6E+uS3qESzBqKWCaOsogB9LY2xuJo0BRNnlbYM4NZHeR1vdOO4ymnockcar+eMF2bhd5AQ
tj1ay1FND+wl+tFPjXmzCHzvtlifGSR5Fx0G3cwI5CQMACn+CFkRVBkZxFYJ4HFg25yZgAOSWv1o
b9od+osFq/jUvYeNa5e9otNg4N870FOvH3fmCShaGuzEWJto3gI7KioqEueHms74yuoKahzHIE0k
sKFz/6YXYQpQaMnEIOY4XpwgBQJOA+LF+FcbUFKvK8n8NweyWwZSH4HSJAqcaHdYHx+acfs4/Ycy
IGKKfKjZPofXIf5XScozZYXIK6uaPvWCestrMdn07B60N+VWEyotD5chSdgESWJ57oi1LTL4bHn4
c834StA7XZqRjHtO31N6iKg1mS+KN3p+a3p0/Xbx+iu0bBrdx33bWsfCCHPl3jPemgLZ4PknxPc4
YHPSpfdno9R7OgwULZNpPrT3HG7T3c5ZbGAJYW7j8/aop4v0MpNA7Rc0ZSMOExvhg3sBwDehIdL8
ZiDVMTbEKzsuvjwW+lIWT+R6EkDkwRK02SjR5v6INOSJG8EDF/gpKy25pgMGIsZyvvKNdmHPmSDc
dneIkhWh2qKd4VLRQeUEHCFIMRTGy8ztsphk0efVyhgWxymy6PiwJ15n28ru0qrwrxDPy6z0pZQp
XwdcPmyPBF6amCbIxupTK0pX/GZS2yhqf2o8PXe8NZVLg0IxMJTWZk83Fy6ukkhsEZ8KSRqMe70h
ezUuDDD06xrMQl8f3d76fjObn2A2hwOTx3CmMwASSDuyUYFmypwyx4CueQAmYQvQTYgpQZuc1EPT
KuRr67+4r8eJcEXF1SDSmKqaxPGGXc30UDrnO7e6tdIdglEAK08DaMTBZJ9eB6mTwfPKAixzpkaQ
t9hioIqlgWG7RNFEzKiPx8HZVRU6x+RTUokia4zNC5jGy5xcGg6orMMXJRnIr2geIcWijaQ7N6zo
bagX7qqELKNMptQE26d81wUYGAxXNZivAYCQ8POU0olqelcb8gXdHOSU+4SffRsAeeMCwxBkORPv
C3AfAnSMpIiAG6YhdBzcFRBPoUX8KfRPRV8jFNIEbImpPsxB6jrHGk7SzfdDzJlAHbxCXqMZ6l30
DrCg9hVxt/Q9ChSGNyjd4uK4qcj7LXj9AWjV/TUIWu1USSDdJ+1zbHRZZ8mKt2vYJRGMn/pRyNlq
b2hOOXm6lWJ9yOQ92KAx2wJQplG54JOU7xgmgS3euKABEbODSEQZ7b4qFtrCiB8yD51JO8DVkBIK
aWe1NoS8FOYnXwnRDl6B7fBqOM417d2wx2ptMkVHPhGuRDvTmTzXTObjMnA5+gflwzVOk5Qd9ZyI
B2kQE2u7QXDfYsdc6bQTxrMM32z6MhZuYJWQWihkDfXZMtoeQ0GoCJY9Qg/gOBhSiuuQKCOn+jyB
eO8dBtq3VEyOS1k+0BTdZ+WFTvU2zkPmUmtNsklxwvDw9cVQRMFXKomCo1Xw2kkBufQPEZponOxr
oEV34fg14n+eisHi9KlCtVCV+8IIlnmm/JU5UlAPI4bRlzAwSUHdradjzZTBMDY0M9rP/tlGQlX2
g7YpLRphg42tUuinA0Fba24t1qC2BeZKu72cB6+FKaikDZKyMPvA4L7LZ4mn5944bOBeWec7Y/P4
PJHV6hZ9wZr6oeTOuig21yK+w2D/rAfJ50YmH0bP9GwKKM0PJ9OnfpI6CiFlkDDDfBQYRWTCULmr
H2hApTFW5+uRs83IZt71HrOmMTW1mYdx9FnYtpZ6+AbwzVF/p+0NRpopvcR74m5yteq/J0W8hyNu
oTMLuqmR6SIyaeEzY+HGzKJVrXc8Yns6LbugtH4tYqNu3mQNYnlrYwVNYZr21aHYWp8J2OcwE0Gy
gVEYj0+uvfam6mjkRTY4k5NfYETAiH4kcHVJC73qNT4Dvx+8sqWW22Q4BoaiHvk1dLR9OiT/e9fu
lMp4554CD/G/oyLaoo1gPEKthW/XD9iNxKy9QHKdneNkxFPffQ3e0vI5VblTtUd3AgOzNkKT5ukN
V7Sdr77Mb6MLP28rIc3aJyJhoHHXgEQTJeaD59KBqw4f9L1ZyGscZsggD45WVvqkJ1GxBPzYqAzN
VCc9ip+WNDAjUrbJqq1bhDO+E5H4L/A/nH69tP41YSwDP4PrPOuOOzYtNP7x1QwE2DCXPXPiaDm6
K7b1C9b+0mumztW8NH5dL8a+cLb/6BLbgO5Oj42v7z+8av4vAzi0r4CFGlclqVh6PLmi6zxolCIY
jseWfpTiFUCazMEgPHLiplAfYoIMAoOILhlsQoc8zFKDpowc/KAdwDsAMEwYeg4zc975Pn8S+eMD
K8OebSWNWvFDjpVbbgg7u8gR1W/0XS0FzVrwwNZzf9IozcRaD0UUiDzgwDijeZSVlILmcYvy1sEA
+RQta638k2D5FIjz3CZY/8N4EXZkmZIRVuH/xVhjnAUrzKDCBa3OphFTUc6M33ODxgYNiIJdm0ND
LLRm281/q4/Xypa+zzwX3w+YeESCDXf+EWxOkmGq98a+J4gjR4ZyHw3MvyvlRlGOiu9hd+4re2q1
BTYpLr9eCeiP6MmHUCoZV+MY6HRHKVgI2NOn1h4AauwxUm8eKBs7Ga7fZN2QpyZCQetkj2DgJc84
C/1+Vn9+qnIWvCGa8e/AlrOc0D3i1MnZrVUV1Nwl5KZ43i/9thVOI/mCYll680i7xyyj66FUNR+I
ZnJVJ+mwvX7jzCL7fiq7XqTzYNuES0OHUH4ZdAfDYfj204rmIYKeXkkp+XrAQp+eUPpU1XMB3Ev6
3FI5aEmuBi0DhEld9kefd5AziheDro0g7iSguP4hpkDEJNUEjO5hydBFz6pyZJh/ZfQCls/7puqL
DBL3ipM3L5CdYWRGQlwh0+U2xOVzoBelkEK1GGbRNaQGMZwrcFxN6hKXt2WRnGIE57mfSMpHAQU2
DXVKnjcLfUX8yBPvDqhgh+DNAodPmUflo7z2hiLQ0hdP6TYFtnVLaR3aGnXYPT2eXrQwcUcw9Uzl
nW76AEakpSCTwxr0FJM+sWfLXuuCt4+IMs4qJGzJJagnM8Yq/cSLhv1Bhe+Au1N3Fwd/XYFKyUaX
Wt9TtI5MtHFU3aj2o3KR7eNPLzkGQjonTl4kPxkW/a89NSyuZpYod5q2yeqT13rb1/73i1dgmWqB
XpLOLrltRYLz0C3LQ/YUEwpKKbJtj2rp/7MOqVEVPzWpYA+EQK9Dxsd/sNM+Mfk6hQAZQlmDHcIa
kZKG/iC04m4ri8DRt0fNvG/1ajK5+rnATY1skkQ0sBgPZ+J28fubsDd9Qt1+J7oJlYk2J65ccafD
ovqUXCcvxgIMDOHu23Suf1SHyZU9re9J+NVbHzWBjqX/UC+j28Kb+BLGrCcd0SZC7Dbe5QAryDye
GPFWlIun4+RkyC44WyvnrEoTgVYGGBfNNZHRbvbIRGgV7/U4O6990XO5XtmdC4J0JP5FtBRWkNG/
2zhTykI4lGy0A1FYKDeAFBadaa8jg+e8tDjxeH7FF8GqjdEFZtsFIQe3xi1il3gGo9V0Mbz8QbSd
CLu+xOiSUAJ8NwoOVt3H6PzBKVZJDWrUG3u6qIFMgRUV62GGmJJ0/ZDbLvH1Tgf5BJB14p2CeeE+
4PrI+Srfr0VTu5lHVnZBlUbQBK0TiV2LxWkHYYQ+fUhNgRB278gay4UOlShY9OeZCMAIrSAH3Wgy
tAO3/A8cnN16Kan3FjODUa8TQAYcE27x6/f8ARg1gLN45ZljC6ZBiyGfmfPLljGXluqMBi4sumUn
Qvcy0zCGoubtE1l92/+Od5eIerZlckHiwmuWNo2OnFu2PJ/FJEZPA/eeLuQFDm5t1zL2ZNPQ40u2
TZOC2M2MTkhwvcnx6tFrSysBVcPglt3bMqdqTN0R6jz4yTI8DxoMc7lBjK110Sgha0MjrvhrzsuV
8tn/EdtlivrL1k80iqrO5ilkc6c4uePzs9cA1G9+jT05ym8Nl4OIL/I7iJyPUI27O2IEKCRD9Y5X
nlt6u4yBfYAKDP9qeu7ZJWAlvgT4SgB8lwvr6vA/Q+s/xmmyldXOpmFi/Uw+pfkvdC2o57LrCNkK
N9Y13p/MroKx6rsoGPYSIOloDKZsrB9No7avdh9LIyT+SWqXm/JWDw8kpCWW2u8YrGD7UFxwLP9+
3gC8jNXOvxBn9cLYSCHCLJ4VzKsqhGathddz/3PEaIDgS+zOGY+7AyLXEksqImNt/nvtDSCwKtFP
Bn/vrd3lMkv9jL7Z+nfzRGR5iSGxuQkPsXN63W6ROLNMIwY6lyeuauBY+lnUb0egghalZdS6gOGE
Ry2nY9w/iGt0j5JJAbCtm8Q3XoztHCrYlu+oCWLimC/vZh4NIs6JcJOXPPdWGAjTLzuFCRizHcuB
GQIokLhFNBia5bMC5L7jFkneiiUCBa8SxCMeZPtHX4kqtg6AvtjNOKDpmkNbjJQG1Cr1ripBKNos
f7NSFU9cMhALYdWddFH+9W4x2kvxT+svIbvwU+0nivTM/ncJui31+L1oWwnrOMw5S1dVTTkLvPlQ
2QAi2RkB2fCR0SxZVITHjKriXkCXs3A33TcL61LXMiQHja/gZkNM0NXc47DJawPTRYqjxj9zdFz+
x/YTOfTXmqBoaV4j+cs8mUKwo/BwGwAakD2bQ6Q/tDGI9H/NkS/BIRbuDZJ687QbldAcZcAefFz7
saZSksHzjGZvwfTRt11RcsEocCGlXam3rF/CK+cAzvcxRQZphZli1t9sj7ZbpFbX3+f5QWmRJOnE
kzijgHl6fCaIvJgQQBqT+upHqVr/d70nVlD0ZIdtl2G8m4K3NyJqYzaRxVM17RrhgbQtjGYhe52v
IWLrIdr+4bzyCxTFvlI7wwS/0kL0v/+NYFCR17onAirAz5xpgNtnlYGrdqSf2wFR4Wwz43ku0qlC
SLOXsjyM6Q0nFBEvFk3WynzRDupVp8XLMY4mdlBa4LUjVb6NJVc8+y53enaL5bwDeLLbmhoEMRuZ
IiiWIZmjHfyX957IaBAmjxHmbTmqdn9V7DPCJUbMFtzIBUpDbVN8QwL3ToKQ3QhvlWTEQwTt2XO3
+izAMxC9qb2IJe519npraqhVLNFDi316/EvnSeUGNhd60hmx3S/FscQXxZMKaWHCOO8qBZ6FGaZo
4Y1mFMT9xyYGMcg60rJiwv82rJcQv/F8Y2Z5+dH0EtwR2WazI2VFLDeUq1grlM9jX3dMRwJt/Ndx
4tfuwMbayhlwLIl2RiGZihDOqnJNzvqc+WYG65+akjSYkEgwBhgPKMN47CdMOH4IeCDXBU9Z57I8
8Om4ZfwLHFy75/lb+gK+bcT4VBHL5OXm6pKEjusM5/E0vuoyVZhJLbcqj43hgN6DQs5ZA+g3daVh
ZRceKoDBnU/ajSrZBU9GNwU5S6igyW1mux/NMMdMQbmeZM1HVWFlRE8KCCS9ffcvsSoTNKmNyBnv
ANEd1kGXEpifYerDjShSliBjkw+EXRvuTBliH+DHuXRxxrqKsY7gLMm5T4Srrrtvya/ktMpK1XHp
yuhkeSJmMa68pKD44DpVc2qmg/QGvzS9dbmMLABY0mx1RJ7+Asa8wJi7FvZ9ywSbH7WoDMueMvr/
pn4c0VY83KstP+oHM5uoIwrienPDM4KEooSOij/jlFQk15yUXEwYGhhQzxhi3fG9dWgxv5o5Lz4s
7lqrxAN28L8EnqMkiqqGKoj32LiZaM/3uluLVQd5/dl2WBNS9WnBybHKwT0IWTUwZ7oAATUsfMhu
W6tWFKOfev5GnUsTTOPww/46qzMEkqOysnHhRa8ibMVUMYEljssZxsk+lyLPfrjUa/JwJxQRfNSo
Fvc32h2GFwwNjMR9b5DR4WTWOM0xUhcN2zcn69oblJbHVW/ulj3mT8NW0avDnm//FAVGJrf19yMz
C/jCNpNGu+iB2hM2IuRqoL67pkKebBSMsOPKd1MT9tV7kmBjWXOu8pjhuHAknx1NwwvdGd+EzsjU
O+Wdy0z0ONW46bWpaxUBlLuSEr6vhaARzjNEtFZXynf6jUbtnvvp8ek6ReA1EPNKnHdiCzCUgS51
hTisPevPFsR6A6RLoSzX72YUILA4aExhMO94hJQlGg2chlCHl7YymJJhDQhlQ+7ecOSltfnVPj5h
IQvf1Xf8KLx7yH3QKo1nsZttpItAVtJdjQvFhKaffjyUq++BorQC8E9TYDKWtaZstnA/Eaj78Nnc
2fJMM4Ao+Hh7CHFu/kX91jTjjKItWxM2ZLeuP9maFtPuxBHZneLLVHKUETuPg3NawYW4ds1f2Izg
Cm4RRANZOGn1MQCZtrhHpkON/ydxHPmBXNbVp7DGOvbe6jxrzAGtrL5sMzUDLln83mIaX3Sc/o4E
SAYR6e8M9K5DoZ6uD74ojjNEuov+1f+XKqG1fpPkNH13bsWUzk22StxU8Iyi7EqhZME6Xuwk/IhK
OIqUOSKLpRlU1ruBquVrTbiFxwHdUSp7WbNgtOMVIT8Cm9H6Nw/S2Aj4/idId3grNPCpqDKwlt71
Sl+CHPGHUnGPNfeGMT5QqpT6hVpGx6GoLPeI+B6GqoMmEG5tUA3MQKylRlxh2DAiH1tG01v3ANyb
lA27q7z0KDqCSRdjk9z9nqOM5yMuP9/d7ISdmZ89B8JXq41xQdqUuYm2EkZxMJXNyjQxSxCewh+4
0nKosTr/NyDh94Ugsz6HIaR5ZfP9mobXzrNfmNlJgzAVNhfgULDDQsT11TTbE0tx6EHrL7R25FwJ
8ihD5oLfqtemzeA1YzbxZuf8YTZ8+wZD19laPmIvhvqq5SFDAJ7MhGfuErDoWPYoRz8KBAKBnw9I
09V+18S+ArJtDV7r3fSW9gCzt9sxLAQnH2lZlylkdyUsbiFdsQxr6AIocEKLEmynmVUK96emBTt9
ZFqlej1vqRXm1L1kElE37rPoEsCiof358LfgMmf7w5hdbaUoZzZGZrebcKZ1Lx8EAlR4UGN6zEPv
H0RBsRl9nXWcDJOfpH657IOPKWuy1p3n+EkLOt2jN8kcL2F3EPHkX2o5B8f1QSvlwX0ghhjXRbUS
Ft5Dc++mEiy2CbGEPxE2NvGfISNLuLlO4SeuaVwyAd/FLBKvRwhKi3ysKkgED0slg5hMTu1GOSwy
17tkIG6lpGKB6izBEtTZ1UlTyJTcMYibMwMiAshPYdThpmfPjRYRnDP86dF8EjxqdNjmqVXRFIcs
X52YT7xCDBNiSPcKgj7Nz6zHg5T1DoEHtCLjhrW41GtCzdk+/ql+OpvsF7NiXI8bsG1GSMkzsylD
Du1DbcPlCPf4DSowNPrySD2JNBszkdW4HGdVGGyPQA48Du+FZfx9tnO9/XxHu90an4fEMqoutopR
wZhubkjvSAg1wJBHke5xSGUA7+/ac34QV9TRTbJLjx8XieA8rxm7BUJaVSQV0agLAVadzZaosJ8S
JzYKaZTFCCFhPTMow+UwX1zZ1N65GDYXBZ2krEIY01RoKr0KBmxHBi+vIddYXGK/ATP7foZE6jEX
4VXg2m1GQRrVMTqiMv4Dp/PilgjqjjuRgm3RxOQRFaxxrjPuz0aYUQYwHmwGtNkq2yuEIRxr6lUG
gee48QCsJ2HBeu8xIdsSfz6bSupU18t+fpOSfizS/d7p8YWAV6brfI3vvMxOoigrOhv1KYQLFkvJ
Wnq1Xz7LodG2w8oC7df63TsTZzKxX/yh6w5rA/QFXDgTj/43F0qMRYFi5B0MD9+jzmHJ+PHj+rAZ
z0nr8WCmyw1dIISiBRLeqWZxXZE/ob6LWHMSI4F2mcyteXiWX/17QcwDCFao8UGqVefmrrMREl4h
5Ej95Cz0/U1PWqKfPiFEHr5ch0/hmSClxXVFB/0bH4x7EEpjNcRVm3RFFKvnG/OW/63CBjJadPw7
dqIsS3zdUAcDNNh6nOodsPouWhLHV5a6ZrM4+aiMlUyCwt68q9gPIuTRpyU1dhztFG21+DgpHOsv
3bh6zRgW9yZ/wTmCKBugpe7Rg/W5OjntoT1sU7ekpwaYtq+cjOgRS5Pg8zAeu3IPyR2G0glURjL5
rdZL/HQE0B1LbUP6+BPXR02qTkpyTsU7IewBgJvd2XA9FnJHuMyOy/3vMoUEALHEsgilo3ob9zGT
fVfv1ek1yV3zCXayEttUbFNTqNt12rvALyaNAw0au6npBhVT1KSmJmWSlvjbO2NIp4lHiCY7Rg7P
V5yMyRwFAQqGQtqrL1KVa2gPuEOR0220QdiAvSqf5DRFIlfMrPQUm+uPuB0w+UoS08FEn8EePLgk
PVWJzohmd4t4MwqvBNw4mAjU71LXx5KgQfCR1pPoeaFI2F1Jb0faUXB+RQKUggYbBE1c8d1gklZi
fkYaBkX7cpxvsV0L0P17Ce8jMD7RpZLkeUcAq7Zun+WnGjFQ+yp75aPcvXg+6Lb2UCgplngrbtfi
/PwFPevgZZ17AHey4xbyt3FglkZbdr6742RFI2zE4W3PZ74zOBnhVImEkuXv0+wE+NzPg7uTMiox
lrqtXnXCQDPwlUVWs6jHn5vn1A9fecgKciA03ogJmIbywF6yslVfZ9ej94B7LBLki8R5jHB9Quy7
3RsV2vTKC/eZr15cVNHydP6XIWV7IDEnDu7Hj5n3EemjsNvOGetnNNU7Q2UZsZ3ncTXN/u3eF/ym
XLjactYyIzUM3SuMSWfKIDZPLQbTEM5RHTcJDtUQ5Tj+byy0zjo8dwYKmJOO+pA8khGGcZ9mJr8m
sbxY/9PW3dWmvLJ0ZiufBgVWWuS2cGAjx25hyJKVYHcRrloWLrpMi9a8/7hMvJ3yK/djsYBu/La2
c12huuh8PXwq6NqInIA2zAII/8JdVoLujrRgW1rLOOshTsRiH65CHg91AuOaq8LhjZpN5C0NcOnn
FVIJWllpDrkRabqCKvymlqr/9rfVDtXlb/Vj9cNvWl/9w1ni1e9VPU5lLTHcbwoDy7Lj+LTBC+Tl
hMai01jMA2j3tZN0u4OQvJu7MSzllIepinPUA3gkGlVX4CUdTejvnKNGLQdiewZsqr/iQT8Itu38
piBRMUtrFweJyaoPrVDPrWYy+jqKJ4HAlbgphssVaG1fqmF6MKF74q/A8MOuWUI7/8OjJNLSonVM
ikfUHOMLZ8tmwyEkKujJYw72L/c2hPOpkKIZ36H66MUhFDIoNF4T5I75NJ6oePv69bC7t7hzLi+p
C1dOTWDr2GK3/+fB5yjLAdhGvkWXXeWH4LPcyPr55yJvmSax3no6g+OVQRKEEVEPYkcYHCTygxE0
vmRK7QCHON6+IBCisSfrUd5Ub4FfKlT5Rm2CRiY1xPV746K84VZl06d/764r89APe25YHKuPyYyn
NIMx+k0zi1j/950SKE6tCeVAlplb87MZvkRdrK1orzZfU4hfGIxY6vFqGl8KEB1UzzEsc/LjcwGs
VovwHfLmBLL7PuVPQtwFlT9FCqBew4n7yN5aQeG1pTQKFF/QQZwkgOHscAYCjrWdmPA5xPvMyQm2
6WBwQWhqa2461JysAQydZPuM5uWD0h8dkiQLC8kYMpbZOh82LHbtr5tpKwlyyozu28/+1YQQOC0y
Ei2QJcH0xCl0ItT48J0kkWf+cVwXNubBcFW2PWxd8JHsN1e69eeZeVWQxSRRIalJeIucMD8uar0G
UAOCY7XSw0XyRfpqXgxaRVnFpL4CwIbxFc2XPb/wmMQpziZHjMdM3WGw9J1B0Qfcq/bxi/9iIuPq
+QiYrLdWO4mVhvrqpMWhv5Ymcj12smb9F67YfMox2sV0cm4ZavsSZw3alnYKzQMZ5sZDVuUPx8Ut
VSH9OpshKOTXH7CKNkVvFgbewoNiNOeCVczJrHshzcaVgxLdjuq2e90TP8jRrolwOr+czfjq+5in
E+IcxC57GNqzNRnfYpgxgO8fvpHOaauKHnKGfXVLBXHpXYWx50f0kB4jHc6QtzQoEuc8EFCXtxvg
CfD/X7INUzCAMEcziXOlNuB03EmTnGDKbtr6eGhnbK91jgxa8ANwZO4521w14SeVtfrcyG0KvayO
A2glmiwe19bVcyZSFXg/fBKwmQOugCBU55QLN7sRuUs4+7elagOnRxKfOpQaIuaJt3Br99pkfjxp
K6O75sSYo9DF4CxOVoAXJPM4QOQHVFai/o+P5F08l5RV5fdo1S75h5qHbUaVE+hr5eNZLKNtMiyX
j8K1jRZQhpjae8NW0ILcn0mC/Q2yn8yQ6/cCAJkCiXEQlZrKBTOVQftwkuNCjXMj5ODv8VlCOY8D
+AxvvIqT9U1YSeudLTMTvNS6issXBudT3oJz75CE2xw2X3LV3N7k4iD5FQaGO/CIdvsTPe3A37Sj
B+6NbfsQvVUd295ljJfxEcgexSqtqM732VoEhrHaQBkQHBxlaIlRL6MsJHIHmd1GZAvhZ3iaJr+5
juuTZWMAx+9FKgDlEyCMrDNuUnVlfa/3jwSPT2AQQ0FjSDGxHtURiqygnaRVMvxxNpKbgrQWH48B
BkQ58meXRJYIBjVxZyjcro86tdoU0lYCeUN0VMh70JgnwV44DOxlgLc+90XkPENx4VMrdhosgfxl
eTt7ROWEqS1xF7rYoZu+5szV6nlClRdoi32L1HsekktIrNCuc7ScgSe3jMjrF3QmHWqKbP+IsHgQ
THi/rjHpiuPf3G6eLIWZWcdKNJt0tkQHSiQB8RyDkQC7lPUoG60zs5Y7dB9mcqubMQlPvrwt+brm
0QVwEylfiqlXkJ7x8wjpRH7ntj8p8U8sn6YSKLtbzEoBEnSV/hz474D9qsT+rVYM+hnGco6OVr6H
/RAiRVJedYhT7kIhF9Dr5qCuu/KLUrih29LTld5X9jAQmuZpcmpWWRWRN0RCdrzhrj7TfO6BLKQH
RRQOp120Ml55wREoLQpoMpsYO6+E8ieKm5JqOievXsBSc8JOPErNQsNuRFVD9Uws5U4newMuR14y
Rj9DybULzx8QQZnws2kcIagd5Usb7TmA5rMJjIkaDRT7cOhq5XrRZTJSdtLr6j+5LNJTTEbRc/YE
Lglo1nfEczsO4UB1ZLzpa8ftfFafJCadlReiwohguSxhfrCjv4zU0S62rldx/LHoYrnN7edSn0Eq
x3O4IW81/14rtfffeViyHcCYAMhlqS1C7eSuvoEZCBoIDxPNprwtPhTpsm4lRbyRW0pENR2ScjK2
Q9vN5KU8kHwhckPjjqyTNYW/Wz8dGDkrb8SVu5YDEmQHISBMvO+xR2GL9xOUehs3ZSWgMSJ4M7nA
Ng+Dv85PlQiKU/3IQdt8BPNKVLcX/iC4NzhnQkHi5o82l1a8q+jsck4CFQLo8RCnV9vJvbA/TUgo
nCgfB+oCGsiznite9RLDcb55ROszDK6E9uC4vzw2WXprJYFivGF659kcdKAfZxVbbyZlNicrvYIE
pRJp/KviFd0GU5i8MBSsNz3Sxy4XJ1ncc+fqrbODfH1rlF1s0/NQ+/t0U+IX16T1yOn/nadUWA78
/1DNf/N/ByGc7c8ji9n+PVTJ9Zmi+F2Vr/JAEkFDETc4bk0GBKa7qS5CRe7If/Ii3nRzgy/x7RnC
2JVmUpuuxD/kmEFPh+v+alsdHFodIu7ysPBnSgcATn2k1JYY7awYGNBZ7XKxoWDOF9Jg3vwENlb1
CwkFq6e2hVQm2RE8Qvjt6LzsyalM3bhVosa6Rf1eyMZs9f0SQ/msxhiJVgnUHZjqKW3r7Dn3TQCo
IewvJfmxiP9PCWIcKYQa9Gg+aoOapMpRrOjjMuoi+Ed9C8ylnqS9BU3MSLwsoORdzMGkixxMETLS
RAc8DgcRF+s/pM5JZBWp6IXCSKLbq4k4y0Sm38VJCr8GDo4b1XxHDs6doxwy+YpEoB9khndNxESY
G8Pcb3liMiSNXGBmoSwBkfe2LsizwjpfMBmRgEnAWlnMZiMOd9vbDmR6KFN5W3/Omvg81n5zd4gU
h/TtBOgT2E2qSCLGewNkBUDwoojsloeBVk0MOlfIesHsrMSdBQKWliI9yn/c87DWsv6D8Drn1J0o
rRd6+1dSuHukq6MZW3NKL/yj7njXUfIUkvsXZfFwfPwEfrkDbatEcr0V17WykJ+EwosATEh1jI3j
3DQj6JgMchNf9v9yto0pTN/TOapzi9etBHq/Wox/EMYqF3Fd4JWuLOy1y/pigpHYVUVx4YXM04mY
3oUOs6WWa5fAXykX9loOD9utRCV83WOfdfKe8WaNbhVt+nFkNpxkAEhXkwJ5vinv156xxlM4kKoU
Gls3ORMJnlr9EOeBsj51HPGciMIzMEW7j6YCEXfOkGlg8f4E5Ftd/KnRIlOj4X+8oXcTkoz3uK9w
hXPbBsMguAs/GN40ZJ0zhqLfqt6wF1xgVMilvFHcjvr18J8D1wscX+/PnQM12DW3i2Ur39td+DnX
929EGcrDnKlfylzgZJ276/HugFoVHp1YO01qzFuXu/xRephw1E9G53p1fZAcHavZrUh6hndfr1h1
vWLp95cgrITqUf02V/2dSzY/vgRdF0DpAEN3igpJilBB/8Zi951lZUk8usFVp4O7QbDzIUMKfx2Z
1cGvv8b7toKmlalFal5Zj9Bm4P6f1Ap3qQVCrhr4ACFVo2ouazBloxJpNUTZWEUmpVGlnvds9Dq6
sEtQ03MT0CBP3qDhb1gGDpei/PI1m5UWy/gT9SGcwy4E0xGWdB2OtXsB3iCHFsrNmlEbAkn+IFpJ
pO8TFIeUShoJD2WtAt/eirMvfAxlSanjU+huzkjQixecH2KHgZct5knVdig+96BiWG7vU0kuuYK3
EIPasQ9wj+o+gierUYvkFJg7x7++qveRH5I9Mb0lfEs1O6j9E1aYBXhjSQkG/n4TNVC6KVmc8jlx
lnPT96TgBav5o8qoeQuC3J7FCl+mO3TZWrs12t0W5Us/P+fN4jqsaeczt2YxQ+UfmwtSHbru5SHA
l9mXDsuVpvEvpZieRn+6dbzHImTexKFV7LWLWuPvDyHLXmI0NGfK3+wMNZPSZdphemPptT/uI0DY
Hpw0dOmWDqTZteIFKfmC8vNAB6iT7hQgCxK6+4IFvgZ3A15nhbkKY/ydIb1J12hDdmLEPJRmhq3+
94yuA2WTUVMMXIk+6LcoAQTqg0b2BRSApgjBzLSFBqAx4p4++9S4bJ4a5ortKHdREwKiebClMVa3
N+aoHtn1fP1+3Zr/3LsMbck5gfFtrnIyB5229AznYlqe/X5xLNSR0wPTuNuhDRocS7GaJ0ckotX9
ZoZFIODqyYQCnn3Q1EJgYT+dBQRqkAdogCV/eK+PdLmQAuOuD4qe71Un2gLFcdJcz4Xy4aqgYlwf
gPR4DL7GBsTq6iOEsebBTZ/0h+2vzzDDeRLUsM/dpsHEx07NWslaNdf79Z5sTU+583cgVIbWMv2h
80vaUHJjMoIDANVIhGwpUKmJaRsEstoZ4tewJh68nDb3r9MR7IVTZ8LI+EjDugHZqDb+B61Aguv6
QFWp+6Usha4AFu2tG4ooxY7sLGMYvGeuI/3hUr5Rtp2WvvTjfLvxisArYsQHFH89JQqr7bGfuNoN
5AcfTbu7SHKyUYzv/p5mPVZxH13CHXyvoM7pA986NU6SoKMyxc5mPzmeJNCoTgt7n7mHeqKHJuV6
YGME01Yv7mFTOyEbiqRR+1/UvGty1KkQGCgMbe1FoGAlu6pbKbLwAC5aMfsHZZFqzAopl/6HhyZG
T5RbHUP7W9vIbqE1lxfUFetDlm6GfBvn41FQ/1voIBdmXb+dRqe0IkC75uxqySd2+P/jJkbgVr1n
xYPj5jU8yXCe7ApIu8vUFrcBC9F8uxeaJCAfV7CmFLBhB3OCqq9sl7x8cOiaaZ7d3vSnFgCSkQDm
eev3NOh7tR1kakIT63h0kDnvOuX7MYgLp0eJlhf9PcXfdSmnIXpukJs/fVabPCDPa6OHp3T0leui
2dhJn4JOfvaUnEZCcwSMyw02PlugtdKFNcNsq4Veqdlusb06ZqLsbFJtC1Jy+dLscYMEMv0xexK5
sEx5gcp/tgdHO3/1uC79AmAnA386JIvHD+Z3H5eiStnv69PcRYfDytWlHvcrUV6daJR0tH4yEyV3
0xJH9GUZfVWwJbTfQcPfQZc5VCQ3tKe47aYh1es3y2rNNW/gPV6IEUP9EunXuXHw67FXvbNO3Ud0
BnjvrTyhgbrVtmbtirr0+Yf0useFZbBPY6ccRuxdJIysPGDEsUoD78ggrcQXlCrYmLbVNdVWbhby
DSulPI29/FjYNc6m9ZgT9oDt1HK2VDAfZQxniZgA/RsMy8tBmX9BsHFIxfyd65p+deBXPhW+HY0g
qE1GD+olmaffXaQ5GSP+Bw/o3WwpW4Im79hrc68rqV2fVGxginwCPoj8vwu2jk4NbdJCh+kQQrNH
2eHq9qKJtXezKgx/gyl960L021JHwLOVaXUmF3p8IXkW6KzUNT9jxJD0kkCzzXeJW1JdjEVq+MDs
0AQlFJD3sFjkOjBCW4ZgAMvcZyxw/r+0MpNJ7ZyKIvB1Tldp2zGLk/ZvZXtbV5ToiHdM1B9EfB1R
J+lOobookXm6h94KUweFoZAxNzr9TvkTpLDJxgBRIxiO7lCyi9ey+L2E9HueF0FX291XM2ZljObb
hwSo9g0r2s34F7PQxnuA/PNWNCmSUkveA88fbIz6ET8XMd+4nAJZn6gP3BRZiUKn87O/ChUdL7Mu
L5dW2g52wooONJxNxgjRKTSlGAemfqCwWwad4a7W3vX9hHKHOmJjjzsPJujVtVTU0ybIuSPXbZRU
NQ0KUiO/5GiVGktnVzaGV9bZkyhcNwzvTXM8N5ZJJnagHKPwoLSvPjj1efS788g2lYh8C0DYCN0e
u+MFEm299vFpz9DcKy4sO2wo/g8Ou/+fMz/vR2jycj7WidsZneib1cN+1tk/UmFuq6/Si2En0vFp
FSyFWzp55SwBD/TNsDoEXVjAOwAfbhWXR6W9qRLgo8ikmfkSpkcfkX1bew8GnALqUyPwDzfl7HX6
ekq4fvJRfzkyXeoVqYZUu82HQWgHriH2WXEwQFKMP4q6G3j7h020cTld9Xo4VOadXa+EIqFY+qSr
HVLMQKC0Zn1tz1JA+UomDpzoLeGgpqZV04ex+q/BrBO850EZ8hHAY9eS/jcsh0sZc2LAlAcd2pxg
yy7knDuoULTo4c4vMqJ7HbY4Xci+nWv3x3dBHRUYx1qzRTx2RgcVWNM1mGmSgNz0yC54rW6/DARx
JyuyVz45tCLW4RbYT2eFcp/iuwoc/7T6cIB49IfPTj8KOEiiDlI0FKXEv1/SJezJP+wMao9++UxX
gckiEGZJg/9uXb9ly5a3MYgIXGYe+eyKFPU1Gh6l0atE5d9AhQntLpVMOfubFyy6/xURLvcYorOg
LSjDqNZ6vr2pm+BdSegONX7XFcIL0iMrubBRE9bWYXy9mj/KUH+D64Ra5HetVR0rrTLZKj/dmBmR
JHAuF1kACc3eoiGJzw5dElmUUyUeR0HT9Fp4AZYvJUP1/G5ppDjzxOhTB/BO8s8oX9qXbQHeaP2Q
Kw/JEXk8MRC/nBHJdXn1AP8t2CeYtdLeWum3fcjMC9XssVTHe2ou/O3UEuhyutQ3NedornkImE2X
CQn1KjUMQJFc8pt9UES91FLGSn9g52rJyfUf+zAyaF99Q+XcUtThs0akA5TgZLGNN8YxQrv6QMm6
29MqFmSZOmmUV9JSeSRIM+tbBpihIOivFw5jn6ZuabGzz9bhjmno7zmOqk2HCFK0sYYzYQCa2U5i
Ykza1C8GNRc70SSUMQiRYHcWVGpIQDVygn+0d/EEm7/sniwuCLckq7zzCpEvaLKm4FzLNK+31M/C
t5PtWuaDS6EOG+EqE4DzbqgkyeX/RoWHT+2ernW5Ixk9QEfXxp3KL9YZhv4IfSwl7p8nfiXnPc+H
Bw4BKR7L+v9WTR/Q/lVIrl+4wyDBqSu1EtWbupiU1s1uTEDw0iZVmhD0A5UbzEnnsmOv/8kGWFnF
mC7npoT/1CeFbHGSIT4mLYvfvU/wKjev2jwqlXHrkn4sqRUfxlXsHK6c2VPpmSwZ3vy2GHOc1Xqg
DTst7BpLgsyjFxlhSzPr8Jow3vXYo0k/oQTXqn6gJdVVkBDuhYaNpzHk8LYmMGvKsbewUdWr7a4s
UGeSArWy6+fwdUEGlgxUXSEzY+P2Es3QSA7n40SN7uRmxOTVWvFSduU8kcCfTXgTQxFLIkeGz3tZ
yjlQoeYBDipSQD/uEEgFDb987YlTDpBaK3q3VmsoFgkcaVXVI+UZBfkGyLPZCTDC3kjJmGL/AhYP
H0su+dKmMJt+KK9wQmr8BOm2ebQtqat2cVwkdmG2G4OIcoUSngYjJjqfOXWOX9A/4u3tXBrG7L1N
P9lK50sz6qnwzUTaTUrxG4ziJ6lUK1yZD3LZ+lCivgQttW264/2mEZTNsRtNWTwLoKTaZEeTw098
se4Kjhnc/sFAbm0ZdOLai+78tbuSMPQncUa32BBJAd+24Ybv06EsEu/pQlA6I05OcwrDtEtVxO9a
EijD0pOxCgL7t7ApAXYW7pq5pH2Ek9Mda7UXTaNIpTvLhWmiE2hAfzeYuzPUXlB7CImHRVqptcKY
j19TqwIrfyTXRuBPg96UN0DIqRdFgGeScoTZzswFPfRTGBRDY7gtV2qyKTMNqWIDutlKaA39wvD4
MrFewVJ9znNyWnvORza/z0K3/S8MFmdhUxosXqW0fMqutRsTJNZbdH7w5uB1gP+789ntN72rrTaP
JbQCbk2Lde8Vmn1anATIHK6VB/ctntUmqCKyDXC8hm2iTXNOoCa99Z2vDjvAYFc9n6W3PGCICBxs
KX9gBvv30rCRjhLg9aRlTFnEr8YfMRkccprD/vA5OO+1fkt7z8I06d0OH7FtNxqkwVZiaq4bHP0Z
xKhtxfsFctgmjRDt8a6WXOOAHzyaneZXMNHiGT1aGpMOmQF49tZQ1mos5Hv7b/34TXtkAbX5462D
kHFoRUsiBZFkGmmFpee33W1I0rDTd+9SCcWD+rEia562bJRHmjEiedej/JfeTc2tFV4RNaFWkBAa
5KAIHGOOkzDKgRTizQpYwEkg756C+Gb4G62pU2IBXdcdummvBw1ul5DEcX31hIFduZuvVJfp0Lle
zbZF2NMfdFLdId4VHYi0uajH00mo8M1YRfkjuT6Y6hBTHs8EPPkTSNgqiws7hR4cGFqDF2Ks3Lrl
2NTHYhZ79/ckQEjhrl6EgwRYCpzA9MS3pCWtzRb1UDEzYHW/WCDdpLvDIYx0GJiYwPCnm2GmRdid
3kEGBslzYWFBNxhn+PJMUgsN/9mr4/ZQkM0emKXtsTUKLoI4HA2tAlmcQtnicbv7SHDopjz3jHmk
Rhn930hQoNpG6lVxSuL1gMY2pauIBX005KGQRXqcFA2OaT2FlFG4T3LWNBZzUBAaimLMrhGOZaPM
BkYorG2gJoU6DH9IY57yUBkLhzsYXGAf6JC6MG0CiMOYg8eY6OmZ3oiVfBxg7+xhirNzoeLW6Nj7
KVtlZvVYEI4XM3F9Xq6qZEgNY5su6MjEGEUYZosw3qFvu/ur+A9RmJM9CdZNYgOjZ36oF/nKBE7e
KUnHhbSxqGuYqvB0O/e5U+lAaiRIhNAOv6x5LgmSgYN6xjFcYZ5AiyZ221FHH4/ati27XLlfUjvI
MTQJQ/thNQme/1AuuIIIxgwulH6ACg6/Kj99Nb8hzpG6cHk1+j7St99VOPhbi2gYrwiilbsAYQ9S
6t6OKwiLqFrEd2S1XcTxFuhlp68kYcxn/SgBvXp2YWzBbLH+6mAP7FcONZsr2cmk8DBQtedzvId4
+ZxbQR5xscay9+DQSHKFIm/4RI91694M1vZUAy34wew+eelcOTHtB6YiTHtUHZbfbQIIARDeNmrX
BVIES9cmGcmOPxnyOqu/WFrsXFYLYDFoxJvXgdnz+l1dPE2GDCK9j/TrsPvHqCpeLPSFRgL7+StC
j+zv+2NOtbdg+XTS930UuZX/szyWjS9HPRhv+VrlKtM2yCaIS367GDadDCR5EZOFEUKl7s+cE+L3
NcevCURg/rxZoQSUV2N5SCZg/M3KRxBiEebYVL6Lt557AEnZGDlILWtioexlRwuU8mfKsy0ate/q
brTfll/KJrHPhbhH2wFkXZFsj+nG0bFFg5z5U+wqAdVHIC05kPUpVzTqJiosXVE5KH7rFpMO6t9x
mitqgWQnajy2w3BY9vAhD6sjbS/xiCk8041fXuNHJ8kOOYIJ5Q98rfbwK33ORrxeRiE6Lmugon6b
cfrHMe31v3cQnhYyP8yCpa9TiWbWmGw0yWfWiOoPAOTlDCEy8fccP5rB5a7jZvVUaRtqDs9BOg1U
GHmsc8qZw4Gq3kSw13bHQf57lzBdrd4Du6Z3RPHO28LFxOw3SU8W21DeO03caNeZ+Ol3z+4rpU38
W/8ap3E3wnILlu4tscRaGEjzQAHfUitAqFNk6pr6i2+oHImAEAFWBHJDqK6j04rYp5KAiFbJ5+N+
Jqkl5ZY/KkJOvGwIqt7IAHCnNhMyffiJQLtDoOtVFtbNM+dJRdgdHK9Zo0eCDbdiVjkx/9Pa0K6i
ySNIUimh/rQW4BtGucxqOwcJVxagp5TFco99RCrtN6giZIfweps0HTPTbs+McEDFs3ngS5vU5dI7
ZNKcYu6I3CkxLnJDyGlIWe8GVUIXfwpsxkMpvMPwpRjBvwVyrL3AIhfvT1+rQyCwqWSjVNEHr+Uh
9jg5N0rZqhhYC6CnrNrd7+yZZzHfb2K+cklIcpWtkEn5QlQjgmNKGgAqIJYnSxLx8EaSYC/611a+
7NYA2UkNtG54L7IKJwAM7GSRx/oN2LD/vrJnYqfiH1oBzE5fETEt+de0aknRxQ2HSGSyWIABNQmZ
BdHdXHJAJ3m6DKvPGSofr305EfZXJThreE/YgbxNqy6C2D5vlLBBEIUfwGPjXnmyVFdWXzkxwpSD
ExCY4stM4TXhoc/OuV9HSyKTiTrqub6NtRn5JR4axGP2iCkLThf6Orca6Vql3Y/6+RiwFtn5+4Mk
fhnHL0tTu0mWWPg3KZg9S7AXfeW7TaAOOpdpzdmQSyy5PxfYVArginl4Om5+p13wnFMG9y04t4ij
bKS0NJczrl4QNCxRAv4Duxr6d0pJ0t7jelc3Vn9hNbvU6dEF1Wb2xtu6LzunNmoh/VFvhQhCToqh
A/qECgABCcQb5r+oA6+BZYc5Qr7mUEplPIRopKoruCR+c1lghdPnezrXx7fBd3l7RF1+zCXKMO7l
QkbYp8caSFi9bcmtLSjFw6ouHisFH2pcUFUhm7AbIoudyJjElplO9seGWHqouC95AO79klUklWFO
ceyRY7t39gK6NWfVjV3bFdQKuwIRPCM6p88PpxXRULhy0k2WFHzcuXSlWj6EK/NoRPEx1oB+Vu02
R6JeRE/MLbjMzhYJbN2QvOXiQ8V+9eK/qL7P/uM33OyaMVUHzeBr3ZtoNsLdIvtWziluWx+1x3bW
fakS53B7T+GZAu8TVjpqyVC9ohlke4b8gfJ9patqPhDxMS+pv0/HFDSqBmMllJ2xkv/g5Ub8tdlu
ny17HSWGOa2yaoBRfvZPiVYwR+eCS30Q3MV68ity2VuaM7uAyghJVZfI0BXwiyLsVrepI/QpgqxS
4lqbN8YXHrTpYCfzdUXePKC/8ZfmtqsKweIh5YyWxwXLJ4OvjP12kZBI4jwZBJxrnxBUOMPZ6uoR
n/7AL0ACPe8MXW+eVlEt3iIRRsDQicsdoeW/RanGhPTMuOHr6A3s2E7Ho/wEL9fYvMhjJ1r8b6A/
w1RexoTlQVZjOnNoshiMWnQ3wHgJQbL2u2WDTU0jwm6RptBUB6n+dL8rGqhn1DoJYvkXadLMvSa+
gmtA+rLkcfo+DtCWfJcb9WTH6Nj/8clfs9E0hfrx7NPESQPqVNzeT01ckUhMWrGR8Fd/KWgdzzgL
gZcMuSzLoRMu602MSoHgNg7fHg/KHWptJymI4WqWPeJ0HRu35sP5hibNKZJtd7EUhlywq6KpQRs0
Re5iuAut0/PILVG5s9IxQTHwAUkg7fyQMmPlgYNnJFKiaXL8JhVDBsnGApU8cv2nnB/QYdTE9uT1
Mfa5yDFF9EISrOe3xjne7V8vRo4Y41GM/U7f4DKIDlYpSe8/eYT2DDdkeq/LKbXZBDqgjMntIJ+8
bZ8p9ibW+ozW8tTMQVwembL2jQQvyMaf2vz+QxxcK7KDv9CsD/7c9uZpPVZ1EHu26NBTfkbPk2fX
EyUlGb89NtXDoBOIDjr43jXGp3sIwWN+8b91cW9yIQs8CNPyCu6FDu4vFMusNT4+EC1zuATV2T8P
FTE9IM/ApCABjGYefOLT00m2GFwCJUrNN6d7L7ySoB68U6az9V8FkLWJZPLD5AddUNUtbtkC5+0F
jrjDPebNFvsTGslI9aUpr0rZ8C0vJxVGvWM1EO2drQlZvV+kypQGx8WtTnFuJjkdHXR+P9ZZIOep
EWIkWnZCfApuftSJMTdXP6hGQKWTZRk7Ch4o9o7hKl5VU6cTgEtx0KZ06sY7iPIR0Gn+ksaG2tb9
G6LqYqb+InT4PGv5WdRtqGFGEg2+4eOaZRE1HczYn64Adxog8iy6hHrM2Bs7lrT37xbE+2VLAgI5
Jhq59xUS1cm5gfhMt2Savg1zQ/bLx7hZx5xftBesyc7qKEwhB/cos25U96CBqQl6BLf6BTyMHKQH
hPwXfe8iIMLFyHqx8o1dG4WhPu3OUm3Rt50JAzBKmjxp+JOsZIbhOuWK92omqv+/AVMdQCmVsQrp
UokEegobXzQSrM0UmUH4ERZVl1H4x0spKsVEnPZl03NHGf1WGHXKu4QYjLBCTv4FRDlnedcvLGdp
z28WD0g+I33mw7URYFlVlOsmduBDbrHltBA+oZTDTjqVpss5+0gSo9IVfCRnn7ohmbIsYK4+x8LW
5XNaBcYubczfhAW7eD8QycW/NDyJ8vGvVtUxQqRYmrVczPnLpwxBOsoh6okZbclP/zvOQHx/ulBM
p/KgCB/wfFkXT9lyFsmvHuNAyZFH/hFwReLPredOLmM4t//RmpL75OvaZgIZCM36RKfOfPSToj4i
43k6gvTNpzgNU1kwdf7uC3Sar0lTmKqdThznxvMG+qgejN/jvkuy7QHM1oX9iohP3ZD40M2o9txh
Bj1tjf3j5jNqMz5Eg5eb/N6g1fvNsO9WyuY0TmBcxV5ADfATu6MSKalnQh5P3jMfz1XLdVCcSATR
qScc5fQ09eckUHkejZnFPFle6ENneN9D8jdeO99sdE2e5Z6qgP7xGoXxJCb1YAZ7CWS1rPzSM3lm
wE8r7Eadsijaj33mWoCDeXdplqO62cHZXA11/ck+Sbv0F68ZkDe1qv0hA4oA06GrzjSkzQn93VG4
cKKDU6ebPEoY8NQLFVNMiIONkXQmgTdpJT3qPblOBNpcik2rc6/HdXmA99UdhA/9vUiaYypc7WCc
bWvj+1XJCyAiQM55MSIKF4KNxd8UAmHl3PoMZnhlsSOMApqaDGSeL7oOBEj7nj7GCX0MI1NO9byz
ZOCjDUQf2cKPBHW55/iKJi+JCXu4ZAwcnvkTwEhXHjBnM9ndpYmPbbBAbYsANbMNFaG9kxGy2pE5
XjC2Lxa50iil3NveJzU/RDCmB5klFZvlBddDGBHrpLNj8Sxtj7ajaQ2NtPCUl5QV3pWME3rv88Sj
CCzCsvzDUmY5fFvHu+2DIrTcgU1i3KcCoFaYEBI7GfegExEoq74AG6KUuPjwrAw8RmqFVJ26Tx5I
uJ6VaHzVho9QHqP7ovrbDsSZIemL1hTExfVRJVpFkwsgEUTgEbXO8rl7hw/Pw40vIfqishnAwSJm
iuRKuFpBm6CYGxFduokaNYz1g3E4mJuMDQxNYlX4zUtiu+/KxJUneWPn+ep3QThUipk6Yz8zVEfl
OsMOwDP3LGAB9A2hZAJ7t7lpLGZeH+s1x6hsMvzhV11juGWJR5YdzQzVOhubp2Qkf+2qDIXyO1H8
iqxblRyOKccbbO10XGdbbkcE6cw+JDUlY4CYJpmSNgEPtRwyqKqaCkKnqSUKW+GKNYERppL+hKIr
4AHLyGpEYO5ELjv2s3K9ty7B67raEt+vpcHweGmCn08Z8Z5V//1Z8SaaBPgLlKGUyFahb7BRqJfL
AEujK73Nvk3kT24nm9YcIqpU1W4Cold3Jr2oIX15GK1SRGR2KbHA8dr7ks+YUgfnV6gJ8URxrnIH
DOefepBhxKROJPMSGdFxin3osggAbIrNpI+PnjLcYABdteROrpk93ryNPJU33iNffaXf65epFFPa
MYyBA5aLHzKCHoTWQ9DbOU6afa/qU2V+0Jo2OYsPDaLEHSuPDktMdnLjnswCijRpOcrTZ+I7oYPI
tv4LXkwqhVFlOwoalEae+OTlgKcTHbinDPg3QtkXxNjeZSANZTMCCOVUic6GG/EB9lsPs+JJo3mM
D6AxAh3M+lZYXNJWFNUUoC+0BDwFyvMAp048Te4Rd6L7UElAfLWUUzX9zyZ40JkbecwQ18zS8k1Q
7vRSuLB757fNl8fkV8R57PTq95nQ//JAsJAv4TBsG+VCMD0wrWBU0gEzjm5wOPcSIgpmB8+VTnzU
rMlm7VQWqRSMdFjz7a14keAG31ybP+jLWmakk0wdnXnA4ua83a5ULK0fSieOcHjmxCRClDXlCSN4
uQwu00aBZ9Ta5Vh+boM7bRJZ+wjuiSUhVJSE8tLNxBM4B3c3mApCST/ZcQ6/Sb6F/wk4hFF6Hb9e
aVoloycfSEytdW8BF3hkD/ZM8p4zsJ4lVs9ulPJfS4wFLSzkG3egcnRI1yQk00wrQxVRiLGeThNz
zPhVwGl+6ZXwcpJb+EiOXdiQtjMtdiypsDdlKq8OUwNf3WC+CNny9t1vxSqMIlVpaoQtOLqlBc5P
FuTMsfBEPTOLYNu61xv2mxoAeY6lzzutLWDIuacYUWB+dOAXKBCTq3BPNq+oS1bPL/kv8RG6F36l
PoK3gt7SW4Kr8ACLw/aVbMMxYwUuk1Eq57+bVsgdrDk6ZvhqJKCWohBPkLczmoFOufRLE2tZ1JNl
Mq+tY3FEj+BjQCLND7yH4ILbR8PXL6sRsXQdQ0CIv4HICsvZYwI3BzQ4r+qh3O35q4d5r1q4YXEm
Th3EQesWBS2v82xkyn8o7M98GBjCbV8+CEuJGfV8bnS8SrTE94DfJV/yGqbnx1J0D4ZP4ShTsiVZ
qN44pOMjpS7MDbMVDpN6/c3RJLvTafvSOovaKQjFEIwFpiR8lg/zIkazs2PbJL6iPCBUKg8TsF2I
9a9hpapJNBLrUosl4cWva0L1U/uAUd80VoMuLVYreXB4NRPfMCOwxxhYGA2H7W3V/A7B1NluBE2f
C21q6rUX2jI8STO8sSCNB3gybxEVmRcOWv+sS4tdAZ2ZTJRNE1BMikm0l5ObnN0vZx32geHd8iWd
YkS1l3X9swJ0QSX7rIUHEs+288gISfszR0Mi6XjKrRbLOEVJO57crRMUXJKTpFX29zBVWmvI6/Yo
1IbCrOdgA5fehEUSo7oFjw78pXUgXgAoNjRFcuHuBXifuqdLPkOrPkaasEdRyWkTgl49lO1hTxk4
mRJIp1baFnchzJd3MWVEmDqPrLPj9bm10Nm13E36O2cNAM9iLHV97q8jUS5Ih92v6Mx3Ipgpq+V5
DI6eBLYRmPSTk4b+rgL+IN/wq1uWLQRUGq0ie3YQDzM0aGRTI6KjOzi1CTPkXFQLnxA8jD5lN/l9
+uY6O1CgxyXMGxY6ae43RAZe2WRnQ4Y0qKdf/1bjsFJbGI3wuTmDOcPOh5EOTqZJj+s6wPkpF1Bb
VPRC2+oxSHOi6gEW1p49MB3ZQ9ykxOCiiaZvnz++3Hq5aIyFMTGbVkI7J6uLXLcMIo3y93dNRtpk
sXOw+axekWRzgu38P97GlFhZYK/uA+FY1rqa8W/ZLMARZNz+OnsKEnej2ovNmzF0gvQUxI/+vWeu
GlFYmVl3RQeorwDBudxdavsvTqS8uxll5/hWfz6SGKrcoS6Fl/4DjmzdSnPAOPD6koUQN23+PCKy
Cr05MAXr0apU7bRoWS+iYml85ffT4/XSVXNHseIb1apYmppngneOt6k6mG9IxkCS4z5TLjsSyeN5
+4Lt+/llpAh3I2ZFtrI/H0OOkqDFsnEwmbUx4PryRXLzvE8XSsAjGjO6PlSVdnf+oXuaa+rubD59
LYfrq5LdFU9Bc4BsTz4DzKTXYelzUYKn90htwKB6zOdGRz0pK0R+in8IZ74+bd9pR26mPNT418Az
uAVy3a/tAUj1UQB0sXbcLDbEwUl4rSNZNjdn/ecXrTEWxZQiMRHCnm5MK8ImRO879j0s1D0uBgPH
TX+ifC9BuM9j+XS5uoQA3vuS/gtNeIxOD8En7oGF29/vegbE+il+Fn71qgPDxlEMVe12FstRwmxy
vmBAY8t694wBWtHcQnKetNWC+S1V8AcSkwImPtjLrpX325Eo1DlmyFoLBXDQbYGJGYPQmPgxerLZ
rbXLYAi7CV88QT6CDbbTfNsFMk0Sb+/Tsk6EZK8M+GBGgqgJMQtbPMJh6qpSPcjlFhYtEn1RlPDQ
f6RFqpT28YoJR6/aNkWAZx3MnHoIPoSt8y0dy7AQjRK6qdInwbUkYnClN7WTAQJ6Gi/5AWHovlIG
AGnR4n+QLtqCSlK62RWoAZ8jGPJAS+Ze6225bTtZMHzhJsdEfapOUXhqCmj5Dqe5dA0gxBZ1cdov
lUuzOBgmSg78ofJ8xKJ7gBBF0c4imZ/rge2/0UxJ3qba8WULohAujILio0BIDTjoFMuUA2PW5J8+
ZdHCcZypQeaPfjeFHm4ELeFTSCWwD7na/2p79UAjY2DfL+7FjAyH+zoEPOSO/lANvmXm88XIYYek
jp8laS1mWuallku6fNmS4WsSPBzaRHpKFEbOBxtz71LKFKgRQPqIfOPzH56TUgFXiKTzwJ6tZ6PT
bw6BKIdwLS1knMT/7LM+VWZGLYusq4YQ0S0mRPMlqQxfDOn1CKOiE0tPXJ1XkcbAZoJjSnzJ/WBM
wwRBjTuWLA2irjP3P3YPQAlBYwDg9FjdKh38ERN2bMmTG9RyaTd+NoZkLhzCoWKOme7y8i2JOWLm
Ma7hWLB+aKfpVzwRUhJmQYgkmpO2wKNgq5U5ArKlYONXfR4iRZHY0MUVpMPytCaOvuyFNuYH2HZc
Rf3SaqzqtHPbkL4UeOfbpbsv+9GVWz0PE45CHJ6fJTl3tK9T0EVNgIKMnIHAUh6BS3dgFr+Ut0M5
1/85yRgFWA2mWhM3asJ5nuMRmFLCSZL9ioBQGiohUm/u3WtD6bSzOZqiqmiC2iCoIREiuOS4PcX7
5qHF1D3dRQhdGTXC/rSpLKxe0bZqelmhhXslS8upy4vaywGeErOhj1GJnUN0GHuB099jy0vvf7H/
+/0mtKaC9G8oRumWJn1oHtvwWbwH0x5Un1dGDfsDn5lvqLiK/uyC2HaGExDy34Ia6TQ1AM5t4w+w
IjuMaQLQhpBjf9Yu2++5eEN1q585C1SS2C+LYs/ARaCIidW0csS+eBdsorILvqpXFmlhNWPFeyDj
P545shsaSUhbB2B8F8t/o7WHRsEuflQV1hTw559pl6R58821PLrAyvO4cE+OPiKK5Th1OfYkMS33
x6MlkNP/qHXKvYpXrhifR0x9vDKB/Jr57Hgj+7hg9E3e+Xa/NdF6zd+0lXMZVjgiZmT30/5KeFg1
9RAeu6Sk3nuERz4fZ399+ezBHGUT/5yyoYTpzG6WVkEG1zCA1s+jbgRFNPTUgbQnKDinoUOMECVv
2DRPOoyvlghgfuKID2qRYAc74pCq5spck1VWZzzvBW+IGLTcWctzDmd7Loltc0yCFhJ9G3omjHn/
mbQueJw5WDQfkGLCil4i7DMeI9dSo/dJFDWozl2bOFRcHcuhlTBdjAmpY5IsNqLAfKcJP5diwzd1
D0RYkESjnkJ50uG0lskeQUeabMywTH6iMInRuGv+QqgcHXF3h4DU4SqN2soVTRTKQxx2YZ8vJjYA
qin6GS6LxVQAuDn/+9yvkNbb7B/WZh5hJkTe3PXW9ShWNVD3WuaFm43t9WcINLUQ9qzjywXl/Y/K
VmdWfUi8WKrpFfkq9BLqISbGm30fOgJ1W3hYOrx7SIytr8z4I5lBuc8t0EcB79WzEz2mBZF2Kt8p
/3aS1DzSYeXF5ZZjhJOIUlZU9WH7OOQAViChB1I5v6iEmCXn8NeZU6yrBEpDR7KCIZy/rTnuGxj5
QxO2IS8gLiV0BinwK/HZHiBZ4HDryZGTXNoUGfu5GBGoEXFdlH4CC2kykTytMi2U5QT5/l7NN3sW
PEQYv0rVBN/mdEZhHXoP5YDAx67+DlDh9XG3jBXgsvXnYmQCyA1Cw5t+zvo4oHhXCb5Mu4SyfD+G
wxUHVxC/k23pN7AfNDc6RAO5WEMGO5ciCnDAnJq3Ux7ImRhfz9IATFg9CmsRIjY78k7uYadePZiS
r8WyWvIybrPaSasZJJ954aS9hAPaTGtW3NbdcUZVv7Zwrszv0vi4zHV0lQaD5my3FQrlPaNcNJIJ
5fTYZHZ9mSqZFPMOYJPjcjsCuY1KJm9LoTbDXO9VU8HkZm5DQ/4NLv3o40GviQCswz4ykO9NpT5c
/aL8XjVc2w2dVc/y4R2h7M25dM4TIs8I4IxFsTT0/sXQQS6pMXyJV8oMO0ejofPfe3VRIZNlmeY4
InHIPp/l4vcvHlEku+j0WC7Ram5/WKf094WswaKegJJx1xHSHSXidGZ/tm1OTn5S3KEB7rDgI9V7
eKSXpvd0thRjVCdFLA6sU73i9qpgx/rQVK+YbfnsvogFuTO2/C64oYT0XYVdYL2RlcOwsSGMCjqF
OA+vLo4XChVox9o1QCVFn0/MbFE2OMTz5a5LtADGQ+I9omYpcssuvX9/k+XSfm2xnrNQwHjOHREx
6GDk1b3mgCcifqjNfAVSLOjqhh2URZPrneba08uX8NLM4dQn6hIdVSxgZVq6VIJw+fpXGJMKbsvF
zer8Er2zmHltxObY0bsbzszf3rwsHVl971zrTTNfXgp7sVtumpmVagJBYfCe7jnIGYRbJswacvV/
89zXYOFgjicUiifxHD7/gfwY25NNhDh7mAUIucNvKMhVeTNj9Af4d6Z9E0BU3WwYRupe4GcrdRCJ
2UHOmz0L/qlbP6tXfB0jUz7qOwvInowk5yoogXYNdTkXxiws60W7upIQVncUFcAIUx6oLIb8yvwl
GLjWmcnX5dQ7YelqefQpgUeP0yY8jwR0VSVL6ZX8X9ONy0IAAU2IZYokVfwpj40JMzt2IL2esL8U
w29i4PWFoHqNNvR3MOpHMfS24gmFfpOC9ACFJ/M0tc7GI/0oW+SUE9hVXhDkL39CaYZ/UT5zpc/u
zyCiH4S2ab2b3IkhLZ3HMcmU2zWc/VB3ebvsU+cm1zrnsILcQXGNgQi+iFk90B8KGqOO8l9Qk+Uq
HnDXvyb8vD4wFagL0mBzo/EkotYIGkFE6SgZ42gDeuozghpAD3eSdPZ8c567F1QNunAsOBigFcuh
75PG5AoQtE4zYB0nYigwpDwfrACwHT8NP/5BYO2haRnGYIl0j+JQq1b+28hY8jSmAK77AjhTilkY
VF6C77yTPU+6wsMSgYju10PLKW1wX/xb/1jvlhKZH9H8sWyeIqPR67mmbyu+v4Qi6sphbCuOzccB
SlLm2/OEbnez122TJ8ggbTtEj3DzQ07qe6Iv+zIhD1dij8BzbFLjiyIdvi8wnfytqqWYUgfYeCEh
yEXJzPBf5KWScgqCB2SoY9DpmBo6T9KpErOkTUB9p5f3sbbCV/dSPBWyAxTziklmqwPdtagUoEcP
jcTMEUC9+XsBKfhkv1aV0PllTOOZRl+vpu5XohS+v5zfhkygbM7jH+KaF82TlKL6xO2+Yo483kE5
riMy7Bty2iDDX2a1jL1WE9SEmqoHg5JtwD7cJjyJc59Ir8EHl6dGBSQYGf/Q8I9LdX7sq1mrqvBw
hv9u7RjbC2TsShLS3njaRcNox3/j9N/ycanjmgR7GbaYiB5lPmN925IglMBzPxJ33wqDixyKyqt+
StYyCXV+CwQEvrV5VWHPkLfxp7F6UHfvHNUwxH4WufkQSU4rL8im5/Yhdz+qLPi3tAbtGexjexgw
ozNGpfD5fdIFu/w0y6PlciRS2AwPU1kkGrEuerK3ma4drdqTN+XYsiyHSF3XzeRyf1oMwEV54oo9
au6CcoAW3cE7sv86o8fy5TcUDsi5rM8RB82hBPopPNyEzNrmQ2Ojo91zWYakcaAGsBpNJFRoNLfV
LLPF659AzP8st4r3xDZfOq5s4AD4IyIqvZWXMZoy+8kKHEJMIXyaIAf065mq4px7iX7xJRENTh5l
6CbSGu6MJGLQ9g6xw3K7uebP4wC9A2hl6nJ1sV2YFAA4wSfsKFL8HC75k4CrmEBr8jVrVCYKSd2l
UbNj31piUBIrAO6VRL0ijfZdy32NLKa04xWVIZ7rzT9sNWiatd56diUChMwimNyfL4k9TWvp0kLN
P2gwmBYDPrzzRw54B7lxBLj6Rncyl+nmu2QSMbU/NFO56ezaaitW+9UbJiWY/ny4cVs1Ixpd9WlI
IZErwnZdjWyEptR2dAOJplMio2L9JDCCWVTcPsg0y4N3whIEUW55OByCJJyLYdmYingluvMaEqQJ
jnwPZViyj0mXvIMjn/84u1xoGb0ApazRJDVY3k/QiuuWIyvhV21LFCILrcYpXyQZWHSRacLWJmbP
nHwwDERA/seJjcBLAglEis3GFveTbex4O9QZ0FPVI6gQZw1f7xprs9gRSYTEo6YRyXo8mGMPiHHQ
Rz3G2xRRzZuHcJh5Dw2noCPUUko6qsFRKtLgnfkDX/dY36MQXZTE9HzcboNdhEBnufSjuFC4gq3i
3nEna+cF+wOY9kRNBqlCqzdjR/zfM44COjDIbxXsxv+UTL7yr1jHBjE9JHOLG8c61+AjYxAKyxeM
0vH1Ps7W+/HIusj9hhG+0AphTFMWrb3+wlu+BJEE2IbX2TtEROaVGCj/Anh2HR0m6l5HNaCj0ZzX
CmRfbkG96z7vlsalRaRlTo4XB0ZdEndNOLNvOcNZ/iZ1AUNc7t2xIHqbvFAo3HZz10Io5G9hZBGT
2WnV68jQoliwV21idVzeiEyY3ZZvIwll5gqtyqVa1MLOoZzokU9WScWa8g02cSGMpIGmmEjBbCxm
pURLvMRtY/O1W1PovqTEnyWcwP3Q2iYaHjmBv4vpXwPaMRSzhMIEUOreok9YfSo3Ts8XZIvu4rXP
6qSLr5i7hTFwdpQwPpzteoA8htSoTPnCA+byYYp8nqmwfLrsn+gMyrhq+Utp4x5Rr6hMzwq0oLIw
HHSUULhJ3E1dDFU5+lWQThn13DZ855x2ELLNfLWgB1ydvy8G6sI1M9V2VAHIfyuBCc7lnhOihmNl
r9yoSHboi00RWmlCbu0KK2jgaoIxyVkL3blj6wpTSYi3Gaum+S8QFFwEE4ZFuTJ/YtFXiNSisPff
1gCTI5gdqHnkxgMBsPImd3wnP46RcVnM1YnXxZERK55nkDCgJ2trNVQSjCOqHbedq7tC84VRGykT
3RNIVsrpt5CXhDhojpK5JtSw5JL10wCzpsrLZh4WL3IU/+/cLKGC3dPJQmSKknI+2Uv5usURGkxM
qD7lkpL9mH8zxG00jvBSj1uRXQdDtS8eb/q02hBFRYWkSddjgchoIvoxeqawd5LG2VX7tjo1c3WJ
rfArFgDh1mIJEqp+h8vlqXTlF+rWBHOBWM6ZyBNcO8bka5J2rlqpbApw+WnicfM4VlWiXxjeotYz
ZuQXIhw0OdSdagw6uneR+ni1mByBtY61EmqsKBGhH4nMVBKrxDiLDzwTgKx/g+eVDrt4p/qJjv9I
zA9sQAtyQZD4Hkky3kGdC4q245v2Ur4S6VogOO6oLHumXXB6lGjVJHS0AsNIGLwD9OwUbjs/LJI7
cWhski0Ir14AHixBAGWW+U6slX0Elwx/rd199k6K3EQyEGMxEoztd59ah6CSGQFuAeIAqrbaGKAJ
SjGd2jbGWmXpMC1BLCyd/tbMMCeUD/ZQHHbc3GOWLuz4VKd+QQdry4K/L28LxLlTVr+FSuj/bi2Y
akiZCEyrC9SAsbvO8/gTAiH4niHV4tjOBWeynIC/4f96WpIwLllgI+QJ96VEVwNDodaPi7Qu+ej8
ix57VtBy1YJ9nmzRMaugjxEpEqUbJ+zrvRu96vMsHbcp1Y8aZvQZJDnvbG17z6I0H+x//9IMvdWv
SUCZgJF04goxjoWI549KCctNXF0pI1XCv6Ao1dSROm1PcTPtSZEIp6A71PIkB7mcPMaVrEo4LZ8h
rlsFsS/ke+KUiPHVOMPtfbENjpHbapHMDzOW5SDW4BHIg8Yq+xdVUPwGrj04LXqvObmRvJBON/jS
E4/qV9hDAC4wVFaQKpXX6k2ftxVm7+LzydTqkhiBhZ15cWvePbPzTNVJvAsP5NK81EuRHSHiSc8a
ZtFLshFInaamYT3j0Eq1JwELE0YVH/DqAM54ltwX22TVFXbAuQZDt7nH2DZds5ntlcscCY/W1wEc
g+8hu+2JSeTe8gs0xZxxnIEPeAJFDVz3NglpQ5JmYkBZVOMXV6ZCt2nzYbWSCXHXfbNFTGDZzPW6
w/vO6X7o7eyb1K4qmz8pWkx2Ev8sHrWaDePmhpgjTrnEbabykZ2c4DHjd5BuX4nazUP13YrdkCgB
JUS59PiYuRyAyqwa5KMvSg/jvKOeuNKnUVNzEspF461KngwNzEYTkFDR/nFu/p/EfDjTF3bIW48R
2+Y5O94/+LBMVYNFPIhVW2F91PSLEVUGSRPDrY7bp0QgP4XrnJKmgjVCkKih3UGFkxXm2UobdujW
kUUp8x0o4mvuEgbJwZNjrnyClBrhPUzR0bhO4jvY74l/geat8NjUrdrU91PAZNXgSzSCl7u0861L
PCK+KJ85VHsGKkNwgQvOAVroJ4A3WR81uPtrW4/mfhedM4uuzIjiIOuE1tHHpMS3cUyQkJ5bgbM8
2PpH0XtCdpWHdUIjxzVUoPNfj9+H1pHbPVNjeUwVlXL6EAXx+BUOqSUu9/1glgR0jeqQnoYbhBoL
ZqIbiIkN2MUOw9n9BwYTjzz3nO+dz/e5L32FyD93aZ0bexcKoj9r5gjHS1k6oxlh1QWzU6/fe2Nb
WYHtpfKBObqsgSisfU8qr5Ps04bUZ340h1pvdlexhdvXDRrLOKJJN7AEpybF8Whh/LgFTBiSaHrR
JUz8dM2+h7NXREkLj+UiGUN3+JUklS06pOpc+Ly1Kq7B4BJ7RHi+AIn2EkRG1lgt0Or+OlOx8IKA
1mc3jR+o6nGAZ3gGReJv6HEuFonuLmT9mGN95Cr3jWhv/eE9Zxvd/US76ytfSg1nJV7m+vUQzUlJ
Zrqlh29H/wBXyq0n+r2EGsyQ5iH7tagqGsCKvAGMbl6EoUw6jFe848mGhwKQW7VnZm9Si/EtDre9
ldpa3ctAQb1N/6YkuJgvgMhX0Nf0/Jbpl+W0eKo9Fgxg9xiTRf9h8LeXQgttnRCx2qit8XMlkPl6
PMcVQQlj3BeueSJAywFRLYH23/n3gKjpZQKThPg3CLDkhBHLhtp/NaZgBYT5AtwtveIgrYflC02W
q/RfaVbcLxtd4p5X6AbYGdOgYlsxqA+8bXzH8k/0pVmSENsiFUlZyD/78SyqgqH9rkTwL4Z2woAo
QdnX677yo71XXVjXIbsEFVvWh4VZTvl+wv0MNWbGKZkAbkITB37v6a4eWILFFvoUkjUou3NPlZ7Q
cL4TdsBos2XJJCX0KvuOOnbbsq8Jyju1l2GebQfn2O4Qeqqs+JCGw35j+648gsvaydKvy50xDiuu
3B1ibR3D/4ta+bC76pDuWTN+dZ8XZEjZOWQDOOzpYKOK21kOT14wgu8r+f2tSpwxQL5WAXpsQ4xT
KtHPqtMJIGiOWXu49Vn6JPFuo6FF1FxL/dFTB7OLG5424WVD5dxEIUF/wy+DLrshVV3Y/6oRjeT3
cH6+KUTrLcXCj1XQSm2At6lcIrJEHHdN1tHI4EuEgkCxwWbHqBNZBfGLaf4Y/kWnPMU/fYksULTv
nr2g6zMz0KrhupphCSrupmeG6SHNoWBREhYmH+TLEYu9enIzg7i54ymD8T9z/cMenFAU3Jgb+NS3
sk99teDyllFmytFe41tgpItPqIxcTWyPB2+kX/57LQmEhcKlthM5SztRHfkFLSMHT0vIrn+5oXRW
qYNnC7YNE01iqFom1hhcq77oTiFAvQmQRKE8kYEhnENaWTuxcaCE2IPjGnmVnzvYpq8QlJM0Cccz
cbOQmLtP5ya7S3oNVk42MX1EsPoBjlBUodDlF+WpSE2UjtCPp75t7f/fRiWytVP4QO8nrVTVBcMU
SbW11OuD/pUxB5geE8obXtTc9ovjiG3y3wLNefGWFw062mGjllfLmn5Yba+uofR73L2sJVtWSdRG
ite3nkkf+yxthptPWa/GU7vpxeeFb+FYoyOEf83flfrBlj30Q7hbjeIYO8+QD2OrUAETc6XP2spk
U9mD8a/iAUIJ0i1xOAgLUNwiqktCkXTs3Vmde0Ro4WXW4rIgs3od83EnCbLjrNsayr1YchlWf0sg
WkuzVc9Dos9XqZkK3uq0kKqb/HAOI3eiAU0F6WhuTTyU0U8If/dwgaVH81o1xs+QvG7N8YSfP4KT
gBw/CmOv5zG3m1eBNg0N/7vw0di//r70bWOS60qCc9IMrZ21N/8lq1CHHHvCsfFG23s2ckr/rAzu
4rNegrtver7iU4tYeJRUd16lKAXmnvZnqbCgcej6cyYloUGSghQylxXqPEX8Ijrg3q1M5V4CT7Ge
QK+9wdG8uz0UjcVZnT0+XYaM9qqrI0xOSPvIwXzai4mjNs2w3d7B9LGmG5FHUUGXoouSOEYbGMWK
ylODUC0/ONWQu+HLrMu43v0aE1BI8mWWPaNNB2xwjBnOQfQuRaE45aLtESGEkyqhio0edtmOD9fA
/u/45BQG1cjeiMdukFt9oRhUcyoUnUIdZhGD3ykud5sGTpyzSxFqHAPRmU3YfD+3s/9q0TVsp7U/
GJ50uTx/mwvXe4JAKKmh4ndhGZPZvh1dKfZycfc3vljFtnvl6V1JZdzL7zd01VKxXckv5yMtC214
GaS0i2Xrbaf0/gKq2lwyc2mDP+2/AsTgVj8hPRSH6xjplybqJfu35/D3Pwp4DgjRDuEnni13q9O/
lY6yuNfZjf4bV7072A1m4KQGWPrpynMUl5uKI1lq09+Rz65L0ANzVSJgeoGu/pqacNHwhGzi8nYU
c5OcXaGArM1vP0gE2QJwkipk6Kgn2uf6YkG2yn2v0bH+JaHN1c7yd613al+LdZAgELPTqpxDFh63
JrL/wn5G+HnI/G+69TQlxQDjIE1rISQweyzi8ais7oEn4SthS7eoT95GFaW+Fb1kbOYSUekLKV1t
vT0y9fc/ixiwrMZb2vSnwSedDdopbduSGLbdaRYBC6RGHPcO8SLqnrIAt4cXUQ/ng1UA7i9lwKWJ
1yDugSn5Cf6LICeMRcph8kubnYsYq5ZpQsDkK1qT6h5nFiN8RZ+gvtf5e6R77Y8DmEysICT+v8ta
+Gb+QW85KKqHrxS0tufbTXAIMmYdRWwdbQsufV5TSnOI4NBvVfnGmgKEg6XrSI2CTyh/FH1XcQos
kzQNxohfmhJDAZye3VUOWSfobA7T7EyeaIcosF/6l4FuyTjIaAx1KfDQwVKU/4HCJ7AiUoeU5rHJ
ZPGg2pZ8JNNoW0Vs0G6hlFtLyjhmLxPScJGm+Eqa651xCl4BNBebfz9SqZr9m+21VUFxJ+x7w4aQ
5RjiUX0HQP9pZVkDXMhTEuajIgHthwxmPlWat+I7oV2yL37AXGueiETUm4Q3oDDlowReaVwI2Upc
4yRfsgOgXnGMbTjsjU3tDu4y7e4BsPI7JIYqxuZ8EkXu4Ong5L//Z89564zYtNNn5iuwbez0oP2J
kKRKIh4zro2NZTYq5z9orKBcqa28Lid1L2YKvNdg8hN14EfDT9tBJJY62ZCDuF720mFLtXAbVRdY
El7qaehRXlUTpC2ihx9ynH43oxPzIyR7gujK2bQw45JcZEXNvtLyN65Ka7XacPoVRtP6BCDzEnX+
uQf+MXW/zaLfbRHHhwnML6N25CUf8Y1EsAccAlLaxZsovmNoHwfL0BH/RHifdni9eB6VGXtt0NBW
pobUWpuiUbE4wKZ2yUzbXaTKjs5erkfbsYNgISxRqHfX28ZzgiWLtxvOJ6deE2TKTpaGteK9coEY
tWqgkK+Kn8iybGgmlvRRANEdRF96/eB+62HJ2X9g16tIC0KsbWthi9WQT4Q2giI/+DtHA485xVnz
fST4o6k1owkNY7HjSCWSkPSKSt31QPT7onu8wAP8uqkdRIyXfdqD5+ui20AvUlJKuDmpiVbnJdJO
uI0ZcOavTJ4GKSTeCAsa4fPjxGVy/5FvwzuQidXaReTfEoRSw9IwIbHQ1wK4gT4Okz1duhQGUEPp
j7Fh61SZmoZYdrbMp0vBG1Ccw9PqOwuZ2hZWp8rTvQn52hu+DZpHWwON5YTINH9dmh/7Bd9nWmtu
PCRs8MgKD9QyaZvU4UM5NgSOUsWLWi8LfNqqaBT1wI566IvjHuH0/xeiohxVzNIQnfHB+XRq/MlX
t/1Qo2gBTh6x2QKv7VvE7xGDIv/gOjvJa9+mot2mVB90aBF4s0+/yww+c7xN6XCQY8gvdomAO+F3
1eyQDT/BQzbILzj23iXp8h6QzZ48PD72AtsnoykuXefcxI7QxCE0EJm4ja7WwpPHU72WACvAVYW5
eLmr4qF8gJGL64sYgXrRB2xD9HgQ283u7GNgakTGSsVBIcRc+6lSDDNfvEhq1hzFLUJzfgKCcA56
OdI9PxRC9yb1tx/GfBBC4pmg1ExsMFteL5iuJLZWKpHAh3EAfXl2x48St2piVnbGAIwMHOZ6Mm/f
skDl7OU3Z8v+gkwDhaBjLUkXvw8EnwHHF7RHb7zLtGhNiv5gYyCX3GbXrplOpXNy8SVYCiCjo5VV
+hBD6YU7A9yd/VRhJ+NQvZ6uoaEKgOh69OmojH5FhI9p9tL8oLXN9esyYEwvW8nWjok6mx7njFv1
UuY3ob4aFRStZzodNKw/1dnScFecgoZ4vUM8mZtxipapzDhCqtugJmtlrY+DKsXrKTmr2xzAVLA3
xy6tOyhiPx6t679h18XX/fntUJr3goOnv0hi2HPy06uEQhW1x+lC+Dyi5TIvqLQ3HHQMQpz5GdcM
NNTidpI5+7V1QEisqmlYs2UsV4ffHDI6NuutSSbKRj4K0uNYyjpp2uRwzfVtoJ7Op/gUERTASXox
efMeVw3iZOBGEmCPoi1aq5m99Wlrq3adaDf4nzHNgx8w1m8OIvWFwzfgDJxPnlIC7u57OztIFlm8
AOWa/A/Ob8XDP5WJG6k+JX1D8fsaWITNaxIqEx/ioGC3uayHjRkrliwgmJt5JOK00ogYYIer3D71
B+ORjrD6W3ddiLPYBLVpDFdygQ/pWTUjq12DlG672XO70HyBDiS6YxcIWhi3E2lnVnj0rPmy9TYa
g14LaygaGyCIt1/7HgKN9WeErpy0C2k3hcrqJHrye90oIEfv2OtbJlTDXbwvfplpFL+jMmuNj1jE
R92uxhfsMETNqAdluMyU78+ykPXIDeOsiNtjPvtsm4nDrXMxGakM+7W0aQ3a/NxTxiUDT4c2Bq77
zmiJh4ENA8CUcg+GJF3kzEonATBSDa5NIPuM2FswMBpA0LFUzAuqIGkUcMYzQDV2KbuRmuFnF45I
G/K7VGkGJM2mdSdM+f2JO9MV4VlaQaVWW07+W/OAC7x5GMwLfr1h/10oes9Fej/nj4j3qmYprRSF
berIypreDi2tb6XcAbVwKknUrkJ76r287RQKr09sS2CdTnfZlssVjY8BXT3t4lNl1dKMwIXcS8RG
5aSDKm+JxR++Zvx7ZWauhHfTBkmL/5xDJI8gKPBz6FeVW9uR8OxB8+pUC3c6vqkrbeMExJ5nYosC
cViZqd2pq85+lmRP9TPVp8p2WpyI+1TYxO2EXKN3k5bnFDztkZDY9po4Y85bc7JASCCTd3lr8+PG
kvDgIqUBDrC92/Zzk2nGOC5qJ/mCdH0+4J8NY7ykLfa5L22MrJbridi7QLaxo5G0FkqZ0e0u6nzO
tObYuZ7B7vxMjz4UJQ01c7oRGVAyf5AjWmuuELySmT2QeVZLSGxFgSD4EGumfwKsbGelVTx6dpms
w4hrjnGe4oVaQEaQa3CY5125jm3Qq9VI63Od6I2sWXSamzuQl+tapNjkoJs9F/36/7bCw0N12bnN
uLWgX7zSz+sf8CAk438Cl6e4vQMIeXPUumdm98DNbSSuZkuwb1Awy71KmvCm2g6GsGMqjuVStN4T
W1YI9uuTHC+GXbLYAneF2Kq3VsjWrfWqCxFWKbpxrd5z3PUXDKgUEF/KxV5QwjR8MZgimucSh94H
6tq5pKvGUTMuggEvmgDYnAkHQJTQdbEtER5BxiJDmZGrN9TN16YKdF3I3+jjNLABuLpYa39FlNbE
HiKzrzauJcQILUgLsPkQNjMN2ElSWorZASifxxFcDPrArWxBLN/iY23gP8XJdvtsYOBv7KRvpWdc
IWG7DpGUY/RvmqhJdrQM7Uas1b8jOb8/8HcoGD3xE760e4kW2+Qyvx/2kqLp+Oa/neOCWF1hUQdh
N4i8wo8pMhc/AwQQFthJbIWr40Ev4SO/QI24GRweqGclSPn4Qj0VoppRrlCWgXZXXW9HVg6bhSL4
HVGReW6BS6aWtIbRmmdqxLjmu5I9g+o82p5B40mfVsqOcpE8bmhJ1UCMcJQvveitkwU0fiX8mQry
k6/1VsRFuFHjcM5ESnjQPoKllGb8NcmDw8zcTEgeraL77/fGDZteUtXfGQiWfZUntS4P+LWluVy0
0UO9K4DRHUVYJn0YmzAdMznyfg0aG7jI4Ko7VJ5ZuSQttgZA4OT75LoxYjp1G+A6fcssaL3auWv9
klCDvkqEAMkmpKZwZEY0pIWQjl8PFFqPDNgXIuz4Wj0iiMVdhtz3ZI0S+E9Z0aOpodGjxb+mUaiF
PLDdbI/VpK28rYBDDKpMpY8zegjVxwzu69MSLTTW1z0vBIB31cy1XHZQDH83fPqkhtbPkpOWf98I
Cn1tIyLVBX229KcW+VH5UGX34VKqKqYFGBsIbU6TFbUpOZb8assiWyFcmmnIDU69kkrqG2NBjRf3
9+rLho/lbESXaUFumePEc6Lan9PhlNWYPM74Yd1yb7ZUglBXHCKzwVHFJBGH3dP3qPBAbHYfK/Q1
gPbeUhl+IN3VieukhnF+dBZN0BUvkCscqJG3Ee6MJoinKdDTZpx8/0NBtPNmePTW7Hebm+yYWkxP
LONtsbDphoKGQ4NGazO76QZG1Zi9tvrXSxFXQr7OHm2J2AImkQtEv6HKeW/s3t8NIREW3620HS/G
SxVHYWQqJTI5S56fge2NBRfn/s7Q9WGueagrf8d6qH34+ZW4nW6WWMTYhk2eGuqKgt6p95IMBlYJ
QsYVWPhI/7Nk8zr8y2fvjS7tuZ40kvbskGHhltWGOiv16EIZdiXJUGxQDMRE/4gouKpOi8/8QHwn
Wu8bmAfmeFXO/QYIWTutvPJP05Pjdux31jpDuj1WlGlJyO3+OjGnbuTxTKCOdkdOk9SO6mmyLXOW
j/xDNaSmDAMFoycrXJGLhsLVj8Zb4FYAgJP5hiKQOQKr0kQEz3RGIGlePze5NmpNBtWX8je9KIP9
5nI/LcpL/gvG4FlGFsdK/a7PYdyte/PBIJrYMYoYPQOAc2LV9J3YNCt0TIwg3/wI92itaaIh/D/I
UlB2VGQaZXuCsd3LgXlv4hq4TA7g0i1q8eblOUkrfQ/3raBW0PAi9FOs3QHlL3WjOsxkPYOKGceO
HSv0FmauyUhzQgkbmMtzSg/EjDvT2J2e3+78KUHKXKObaKdyvDKVtsoJsJYfJnR5cCrjawM0Fuef
nqa+OGc1wV0NTjjl4nyJunL5PiOYXYTZe+NzHjQchDQx1P/je8213HWT/pHcqY+o0FV+tnj/FZ41
UVPm6SBKczAggi4BQ7RXE2N7juMPr5jiGNC2tahCtsRiTlBBfgpJTUC54LVG44+LdrzaHe11PDIy
j7nuKcERvpRy5vzgtVoOzAmt/urH7eldoJ9V0EYFEoE56D9mM7Abcdv+CULZGAnMzT6cQSslfqXC
f85tn0g7z3gBQainIX3HLSEqNl43h91+dPQTuFOKvWc723PrNEIR00Pu+Hv3hEPz0XRzUtWsxd/s
PMwkEdRHKHBFNbVgVeQCjlcdL/WZpMxOSkX3q8A1iu6SulR/1sLdSBHfQb1vka3VVoC5SmjUfOXr
jDO3q4ZMbhhuK6POmtuUyeQRZtLgQvJay9e9wa/pw2hVu05+m93R7N/pm0JPURTeniTu7/tPuDAl
uhDHehJ2Q11rtqOtSUxfbMZC6z3MO6hp3KbLYKNhAxTq0pAT6ZEoXq0SvzZiUi3aNMlAYkr20r8K
EYgfZADXramJ2AtxqgC5Nzr0NZvgAKnB6JJL9AyGhKwBNSURib53eukyIanBtkaTX3WRG4s6LG4h
kOUKQT828l180IcEYgUPCQraNRoicpJXkt6RSmXGDf6Um4yKcojcewRgj6h21bMa7RhJUMF6QABG
LHAOVlaD0zVQR56SSjZDVR96Ni+w4rlNzgXEoGKVGS/8Znn69UFaR7Aj6ncsdS+Hj+vIBIQqr2Lt
2SAUJwo4/kV++hee/St/mnJYgnyvz9DdDZVCuJJ1Stv6Z2R9eq0+KisxE1Gymvy2AcCz9tf6XQEd
TGG7lBETqeXXMk6v431uVjMfbtbRB8Xc4a0V/VBJb2rObQw2Y3cOZ8IR/lLit6BIxIbV+tOYqmay
f4wMCAp+r0kxVV1ZhmYTKL7qvEgGUheIsUrgjq9QMt5ewkqGR5Y68Hm3RNNAu/pjtbrTt2rtBHAk
nvtPq6g1V9s3pc7MpDXp2/rajPqM0uwf71EzHpgrZzpXlvH0uDXwcWOS0oc3chK/161qKQd1EiXI
9SgTAHVG+QXcYl1ZtpfsX3/FknGQVbtDJG33zzotzivyhhaFnuIZcEKEWsSgllLU3zQnmBEbvP9V
lXWZcojkOHplwmTjwKfYG7ActKZlNVfLdPIFroWWE5b47QQJEJQliPlB6yr/q+0MJJjbITxrXqUI
s+Nz44nWqMHOrdijDIIs+os3oHiOHjaLNfiL/PLCD4h6H/YM1rhNoflhb/gZa7Bv6qIbiPUcjDoM
bkPkBS5XAzdQ27384B54RJv0skP+5esxxaDfK5qr3YboppR0C0pd69n48ahCUacsJG3OdsLH72KX
2CybWoSDE4TObffx4iViCQZoESf1Iw9hqYLa3iTK0AoadicyXw8ZKgEgvHi+7jMRae3z6dq7VLYY
J79iQWZ9ywcfKDyJ5jtfBeP7cqyfxLNlpv70oDXPJMxJ4sI2vzRNXoJdFL7YJ7LhLq1Yaq4NETbm
X/zaj8XNfr9OmGIcEcxofcVy93MJu6EeL+QiNaXabId5CN87KRMgm5fB1CwLXjbOVe0pU/BQTFGF
nfJcJsGVccvH8A9XjVIiSsqRH4MBIhkW7DjPKSBdDhoTiP4AZIFwNjc7OUqRvjQecax5q87L45kv
7iE3oHj1Gkt7CTKUbBtF7MVFdmGwsX1IyBjJ7f/t1pgljczdPipYV9hEY9KSgQvWHZc2lpUrmp/c
PY83OEYJjqh1ocGX2gJfvMmzLhOHDLvBU3XkJnOo60d/lOREx/qlzrxbBNT1hfiGztKo4L+adBBa
K7uwTzrjE/nw74HigZk1XvkJo33g54BLk9wpEV3ravN5VYAmTTurYkE/1so17oSryjX1OXyfaU7F
rv+933h/sKpt47faxFNuQkH3wx9YuK/JZsiAwgUFofJHZBSd/uIZLqwV4OnwqJ9NCoWh93iNwZoy
eYGufRO37NpSsJgp7kovHTKVcFfyU6F0ykdWBLF6ri7AShY84BzceRlx2V0cjth926bIhFg21COF
2ZjexvJx2AHhSVUvEjFZCaRixt0xLeed2QRKwbFU36wylS7s4IY+mKlACMZVUYg0yx9D5G9NflTL
l0wZTp06P2+cRUn+i+eJiAZn5c6SBIy/BiB+eSpq+GYRTIFeyI/PYCXp0UFL4lgpd7/30/O352ad
MX+v2QsBSW9dUh1JRS5DOE5jEENCJl3eu2Oc4AtBs4J+JZr/NtvetOKrqnkhtbhh7RAnTtlMeTeF
ExJ1CbqDbX2Bbh+gAhVvLq/4UwhEie/Z8cDWFc6BucwmUA7ZGtDK5vyznK3uCW/xToFy4Mj9ZRJc
ysGedQeom022kgfCZeZwMDOy3W+1vwbm8PCAS5r3xiiTvQY5xYw9xH76EG9mEMPc1gn7/1yPQg6q
1rImGCf1dVpRlM0xrx5qoGLRc8vt+bFB6VPuJ9SWlJ4o1D5mNKqjyNdzvX6QX0mMaEFpda1De4/B
jqdqdvv7x6vdZ+5lodKU74ssFutT5uBwhS2kQyMrrSZdW+dN0fHYof49BdRlC7cNNsTiGoytI1Ni
CCsic7dR8bDZS7vP0QPZaqJCa4tRlNqYHsEUWg67PhGFvRImc4YfuNqgV/ukseNF+JyrsSv/a+Ey
jmFC1S1C4JKPAHukXj8JkA8KoCiku85Ja+rTENwt1vPjyw5a80c9wLSF3taXvKQd/oLdO/lnDuzF
S+6qNu0u3ljsrMCKEHLWsVSCagUBavy+z5By7fvVDwLONfEoe3MYGsuDDkSy9Ozig9Sn6CAvg/N9
fs2pKkU4UqkjyzLpIVRyjny8ZS6+K+xcN0pmknIwBjUVuEupG4SPCMYsEq+v7xXs7+IkZTkhc1wg
YUmnk+thIRvuSmoFlF2U1kdZnytFrE3d8KNeKm8wEzejpodplJ7ulZHsexV0uNq/jjflwzDxbXub
YjXld5y9gMoThVHsK+bLI3+SULcE4rUnRCnbW4dP9gecH5Q2pT6i4icrPonNAtowkYNM2hDSipL6
Cx10mori1RDm8zBtq+c/Po1wyvxanQCY+mV4CI2wCEZn5+ze0FN237mDVHo3lPuOy54o7DCe92Vc
u+3TSQlMU5bHWzUP/U95nmps+oPAtEFCWgUllA1keQahZnr1Gsrs4STwXDGADavRoACK4lwGPBvf
3OChnFQjXpcaiH3CSPiwn2Uscb8sC8bYn9Uqs3j8WtR1w8HSGIVDNRDecJtOFmtkguAmxmxEGcpG
q2/7ThX5y1OnkQnHe3fhZdDY4u0Q5awWYKMAuCyPRmdiJ8ko5hRpuA+IXiQqwdTgnfI9KVW2qkKT
KJAVRcVRrlF7WcVLzfOoMC34fW2CyNZUCicYkIk6f2PxuA1AgPNFi6k9HMC67w8/S5jj3sUQj0au
1InOuJXwpvQkOtIIrHIX0fMKJj1VyOypzngL2/CqLSbQPkZQ9AwPS1yM5lp+1mQP6SS0FH0FoqHq
9XB/PIbvI0VNNOqs9OZkUfC89RVBNtGetjKTQeiwqiFernqMTcMv1Mu1YRlF2gXEzhcN2ejoILha
HWpDNAnHdc+k+Hmp3zGgxyEJmR6+K+hgibztz+UoB7pzsDr4KwFb6b/e35FTW6gofzfksbgdJ1S1
GBKjzwERzyERxqURtZa6uXwGDxzRelfqGKJl3VznuKL8vhIsR5jq7nV1z5K3YDilNFr+JpY9Q93w
zntH/LsiQ0eAg1gXJI/ct0mHeTdOPCCPjwb4JSJuHQV6hiJoyh1zuegxoPEM/sMmQVFfvSlIKhLc
+32AL8kMpkI9ls8yrjkFT0GlrSylqdQ1Qp9seWHE6f6pElmL446tO/xd1xcyZlRd5bRXtQQg4yY/
W4FNgUwk/dS5WRHnGNPAP6uxBTYWp+4O6z5JdQvXholvOWkkfo/qBOj1o1JtSSTv4UWvCUrm43YN
9QcsWhNKPlPix/RN8sLb1/g08OK9GcynpWSm+RdETMzZpqrdMr7wyWrgHU+5nHSr3eDQ7pXDbWT+
kman7YehWNzdvG/kJR1QEEOwc+5QjLeAaPdJAhg1MpvhqFaIqnywsZtMGlDh0ORz6Kix3fdl7vVQ
s69J5jI961YYCQaMR0xvLdLmceAYagfMxP8FsoeD16ga4G2Oe7seyJbGQa+ElGuoUlZaRgCd4BRg
uEm464Y01tXzYx0H/P0xf8wHobl8o5A3a+JpxDDDcXtwdqeOZH5Ib1DKwYkkJmeGLv/ufO6XjzXr
TpCpZvyF5yLygvLM0kviTYPcxEkSMiTe7aEmaHMLXQ/duvoaN+eG5rYjTdXadgft/Q+5tISlBo8f
hNoWMwARuR06CE7IFLprZyiKCSoSpVlLrmyPQ4URw6nFqKnLNL0YIscof+Un9ckGJP9RvrIg4L0R
gMUq6OMsTbj0v4MZ4vsjiXk3PUrfAPBdzo+Wla7I8DuvsKrX4dHhGDEJUhB5XPsDX3bA4TvL/6Nk
scIp1/TSmXmWUa4WiCZvE9+PM3XTFf8PFly9+YQ6nktHqbwfcIlIwjgUupHtRldmhKU0R+BHnwlQ
EYlVs8NiX1VDuM3j9JRIHxe//QwbJPgLrjtMa/B2Hblmdwkz1mS7a0IRV7emsCPI8MG64NLWST41
P7Si799YItTKZkp9k+55hx3n3wnNV8Lpgvkk7VCGjf3FsCOAmz4kzk4zcE/9EQDxojTlqlgKh8/u
Xu01wwsZJ+A9TLlUqckPqpf+Un339yqAv1aTpDP6jfDlSGIdMWdSoQrQfV6h65W0sgxncf7BlmJi
8DhsdkwI2QfEdgmDKL7SsOJujU81MchDyweQS29Rtpcyr8ngiIui0nGgjeGZMd0Wd+SgU8UfRo7h
Df7prc2Eu7b5j+Cc7KdTYNRLGUXn4wTR7s1N5IAmuqnMD/cPJ5OiNgpXckk2DJG6/U3cjvZCaaBs
DwtBN/ivRoggyltjJ1xiGdz1ZxzPOqMm8XzyaggbmHUJDp8Hd85UbwbDMVCDN+RjABtj1i0e14s+
IVq0tZeRTPcktiTlcF1W/VkYwCTdGXrdhfFUSUP0745hCqCPVz1U8XmKgYtIZ67GC5DI0TBTxnZF
yN4dee2nYjfEXwRT3p/EXgmm+L3S/SCDPi+Xpv3qj/BZRglgVsd+ZoPFiLVwIwD2d6KhHf2MFr0N
eaZfckgWrEvXXoSSTwUqYI2YkXWpKxmPdR18XDMYXGxwHRbbnilAQTzMv31RITBr0AoUrIhvzYjj
tRTLU6Bp4YDh9OZCKtoe92MKmAOGOg5Gk2s7fpHmgB0W+oZTvcxWxgIYavz4IhepRyJvSBatASe5
qpW9TNdZJ34E5SUjrvbvNbHay5VXZQj4uBRy7Jj/1jjob6eEQZ7IJCuNiQKdoZboTHL2VZYtHlxV
+X/VvpyovOgqsINOdvsWfIOOowFz0iUnWemV3nH8i4lJc/y4c/CkTU5/MBFf109MKw0A94fGvzpg
D+//2PwrOeXCXp8J/dFrVLrG0YFm5kqO7kZ8GKMjlCGzRiZxgT/CkwsRybny1/ayk7Qn6m1h9nyI
qSW7jBELOD9Hr3jhJlmqNVWSHoHmtwKgcDwxsJMQVnxlRQ+7TUwsM31D/BEkDBineidSnUVbuzHZ
UG4P3FXrHNGXF/V8CEWgF3TPpM3bGgjlTnBZRrrX8G8rR3VFx/rhVM7H8e2pueMqKiCMfx2S+UVw
mbT/o575nF34pGVOFm769ofhgp1U9O6TjaQxiFCl79hYwFeGUo4A8H19dl6bXbDSPTodp8aBX8it
/cD1DWzTbxs3D1uJMBs3ePYgLtPN9WWGYutMTYpOSwL4Nv1D1h9NPUDd7YQwIxsTFWSc3wX41DnX
r73peHJKjcJBDbh5wjr8B1x4gv4oQLk6BQqIvxwqn+74LT2ocLrLqZ1nGO5WlXhGTZFEYvuzYXRl
Srbs3/bI3LA/fmm3ZAzZ05STxkdb+DcYeEZPzlp2HtALMLpzkCabs5Bhm16jsJ4w3kYOjeKPvxYE
oMo1Wm4alKrJcRSUF7tlzMqlsqhc/n7vgDxZZPyU7Nt51yvOgsJE9Q/M+TGdWnzKVQi1pKFAHyOr
eHjtP6dP7UdYl7THLnDjNpbg0FQ3CvdqUzPPJqCXtKFZLMiTH1hbkon8NsawnS/EqhaVbPcisCHX
iZwQNvDG7fzeZs1e1XYsGo4gmlupSnupBO1zfMHh0M2JjUEphF4PWS48vW70Fe0rRZ7PX4XRt2Ee
h+xosqPZU6gkN8BMdP0FFso+GRc9Lxu6FKsCKyCOy3D341APRGJycEA4nFv7DmVJICSFNb/O6miy
UFLeHXf7rOQRT7Om2uJJPtCBJlLcnY+Wu9kaBumuHnJ2cKhm23KNuvyQwYQBDBx73dBq3U+Xy82T
WKlK+YuAi4pnfhZcTvC17eXuONSQOYEhKfTK+vwGEE8/Cp3RkwdZmZ6rmsSkTXviMwBQw49sXO6y
fmCbJ01zzgTZp9KdAMXQ8k941/dgIjKtlApz4e+vGWPjiPK12dAq9J9sGAKKIYM48DPu4SsKsyn0
woK+gdBG7QW5GXGa/ZqMsQTvQk0kteFWZlh6d4MFGiUjzfz1q8VQ/DpfyGt2BBg2aI/p01Rk/dEV
4JsRYoRWD+i/6F7UEzpdkpdVptKi4BLk8RqjqPLmiPnVfpran/OjcpKsohVgI3eDWsmPdHfFE5Ow
dI91aV0dX5QUTpHfwPmZId/CohJRS7NUi6WBRIIoS7bZp07cxJbdepGNdxOFfd3MUhFFPryNCdjW
TCurmxHfQXLFZK9RdFNAbjqT7ZbunJNwWlNJgZvzDavttDzrEFWL7cVMDsvLOGPKfM1mkfjkL5w/
ofR2pIEVq+/vg5RHK5W6iE/+KKjiLTl0iHin93pt/1O2r6m8dk2IfPWQfowK3fQ5xDuCClf4za0G
pCmxrao5WPcdRLj/ZRmZsDV7b/roRExqgyvLOCrYFmE2WxQ9cxkFN3VYP1AWl2zdE/nU4f9VvTVF
JQlrc0mM9Rl3PESOholrxRLJiA1b+yAEplfHpWfIV+MKW64J+5qFSngCHJQMlAtkLdfz1AgVn3Bm
1nsM+vHfxpnu02q/CMQndbuv9QRJxbFJrOX/r15CJqWXFmbkKq4zbfhxTPbppW5JYiWANrhKlkxV
abkD7xitu5NXU4pKjv0791XqeKqJEVC0lXSUEtjkg+aWWwEAIYPAvBAQzths6u7K2Eb+KdMSuT8u
4quGeme6yWiooWoyNcen4pmkwmS5Miq9rv+6HKNjaINlyPj7sUCmtkuIZCBMxr9kF3rMCc/KQu/l
1QeHMInFkFhHv5Z2ZYHVrq9l2q5gC/sFQxQJ39vmaSYEoXbaWI6pP9kEIfN29jgjkNhe8DX3CvmJ
K+6CGUbiew/5OrvwxWiWW7opqowkYitwteTQDQeobws8J3lqPRxuEcrBDfufjnBl0niD36BK/suW
n6KDlTSXUzaxv6u8VB/VfS278euOx7vmuPYyif0BCAZ04NhLTEXGSxtRBha2evTurF+77SrUGGyX
GCT2KNPYolHoss7FPOojJuRV5ecVtiiAB7LsUVDEAUPwB2UpE9VodYSlrSO3xaTm1fcI00zPlLD6
aCSn+6C1UUzUe4rBEJG4HTymL4C0fpeYrJifVaz3iYCXJGkbuUa0GQYNqv0w8QqCAullU9bG368Y
cMMywOYCqv4f3mWQu1epeEVkezwiP2GE6zB63IiOf2Ztthz5eQS1JRTbu7vu18Ykgmf7O9xxY8Uc
LoDkE8srzBgQDfXuQVFddjJeea6RlNBEhKQGv7BIiPWh2qsnGS+U8VoPF6BE4wLkqtVgHU7Or7fA
WW/SLR4LlasYa3kJGmtxJBgBy9YlwN+kig+EdCNhVk+V2Js/LE9lzF7M00FQRXXl689JqcUfEhQz
AqMu/xjDRtuIuIC7LeK9wKESezBDg8M9huDXvVOSlDb8oYgrFGlOmSLDWEQeJxJwk1AIsZNf1/0d
qUQkbjhxDRhoG/+r1fWtSZZeq/IAAG/ikTjDutg4+W9KUW5SjMEfzgac/5Fk8X6obFwKoCRbKlv6
pp8bBjT/T5W9gLg1i9gMmREXpdhM2kBOAmqE0L7nHd/XW13p3s9604synkup6kT/qP6uGop3txu/
vmmM2ezPVssfKLVw+5DRPvRUSIslk+cwK1FYpS0WnQSJ/57rAACQCqJQcUQttoxus2Ip1GwE5u6Y
JMymz9EQ742krauVGHU592wnWbSPB+79sEr3F2M5AWm+UdHJa17yXqA4REFMnh3L3Bo5qwY3vbK8
Unt/job2/JJAUL0NZg8ycZhRZqYGJJ3dToIFrkgONBdxvHt5MZS9dxGg3Lkyk4Rl/3C7DmkdB5Yb
GRWgp1jvUe+lM/edUHhJ0lEbCvl73czA/HRSMPIxIk8hVRC9EmUFR/mx6DUxh/W4DqlXbE5j9Kqx
tPoEzAWIWskut2btO545AujixlF+qNswt0N12tGA8NbcMEwtj9w8uGZUw0n7T4utwux1/BcU9tVS
XJEjp/ssO8nkOK2DlGcruOxmGYW433vt/Q9SioRRjeUUotYkSk9ZFTy8Q2yq4HeirEeV4692QVIH
rpzuYb5uE5CGu3v/XfGofJZN9JSwc3l/D1EmQJD0sBtO9lqjP4ONL398LLYA2btQHk3CV5k1DmSB
h+3h5PCaQo1ciQwGUqUIR9/K2MvmBUUkC8nWv+6UBQl2+IJyXHEseC73qfezyPJVYFTcZjz4K0Gd
UPCZHRoJ0Hql6LK1pLbd7oU/CPTY5cegu70Nv2sES8ZiECy50d4pFscYL5kp7Uw6R8egwR5Ont2H
P7Sl+YzfnDG03FNIXWu0ze3ZHCVhfy4cXloXWz3Td5HlBJQOLDW/dZS3vvB+Xt2KAUQ4yvkEhOG1
nk9SSj1VKRq5UipDzNFgzEN3haYnnlSZUIxnbfNlizPi465nqi882s8cOtmBmYI4cAVtkxM8rxxt
kgS4bT9u4y73Bvzi2+w31t+g/IslVxeXVl3RKyUslSASwFU06NgBNp/STfFXueRHG4ffr6Tbd5Ll
VhhnUBEkPXRtQIoHRBS9+xPTcjMj6wS4fKm2DAbc35ybBwFngyZuJ0ywDwhT5BEyT3o4fVD1ZURU
W8zjbtXIzlMWimVj3kgLQCk+BLf+u0onRHcAux+l9Qz9wVlnX2dmCYmYbs40s59/0DXMwV9dCas+
ad3/J6I/NtVmGl5F/1Bc2zJ8BxnrJ5QuRDA8GX0cYg3/NDl8GvZ+fo9qrr/Jg/nB3LnjvbAYzcN2
BcKpxEpWgB/+QDxkERyPzaz4SarLK05DXiI+188Rb6ov1GyD6EbJjaTtGBtLsk0FLkQKLLLiZiyO
Q1jGJvH0guiQ5l2+npHJ84fMSPnkc3cubA7fAvbpL/oqbVq7d7yJJMnzyYCR+N5joRwHQ2iNmTuS
IfUUDtZPX20sHe8WAjdiSPQB3gn/o5RLe4n8SRTZ9hXqbbXms0o62W06E7h1FxSaPbGnmBP8Db0y
gscSJoaF/rPd0zKoimNmctuRnzWt+EaWHSlOubDNhMDC+gXxWP76VTsAhyDRF+DaOa3rxVjxH/ws
TfF1mkLihr4pzYPjwnhkpy8Iu5AlVv4dX4Zxklsv5/ASX2vjDNUh4Wo8Ewy/x6ErN3QJhGjeY4x4
EewFrQFwwXgjofaKgFraTsLTVfJ83ZmNTYMmo6UoZOoH62rh2i9sT6W2wMJMhGHac/xWQCB36stK
4R0eT3rXIeFqw6CkYVFvHdGftnd67OgQ57ieY1O/oDklZRAN8Rj5coiN99hIGanZG6zqFcijFUWu
AnYBhXKmULZKGSgpJBsbV6hlqE7K/z1h+HJ24N3UfwLV/QThlQGfEBvcuVhsh8J1+MzAzj6ff4Wh
5CwgbF+yiHak//r+eBsevQ9Z/FHpDEV/JGR02UbMXdlUwnTt8CH2aworZv2up1j2n5lM5vgKcY9t
X6zMo4Qp2swFEf8TQMNaWRQBAlDah9JMoCsB369oLL8p+EeThzl/Xd8z1AdgaSUYqEkLMtdlSbKp
gZsUybJWedzoOFb2IjWJmgeRZty+g8EzvuRx3FcN9eT7TPPHvqVjjLETR6BI0x+ChVSJtR/MX+2R
SYMA/sQUkR8SV4xB3hcCSLubksahzjevk81uMohRbEgnslKItbpnl61+AICDA7XxQyD3SdsiJp9k
tjoPmuwBB6K2aNQQKEzca/Mh7sqb+0owJGBwaJwqKwBBTmlJiEF4UhJolgl8WkT0/833OB27t3yp
rXMqb6oQTlGQYPykvWxP/ZSSC3l+Bf/Jk5CjKgQPKi6VnOi/IGQ4CZ59xSdv1AVzvZNj6qILki/l
i2KGM0G9dMKLdiox1ex0XkrHxLfsH+6yi8Ys/c/AQO8gQ/aRTdnwxR6t1F8Ods2yj4VBKtsHarhH
9sPXt2TReaEgPyzmp56h7Am9IkGc5VnbU1sN3d0zXgeLSRC9qLrkvlA1jHNGiFKzcNRWBBE+iGG5
CWoXS7Y9bWXAy3UKifnLDHngPSI8+HOSn1CnGsmDIKLC3H/e+P6nP1w+hr2nzG1TSlWIcSJ7/ysl
SXgHNeQwd9Z0fVhXkAgGInptMY2vxbc0aEIXfktFpoCMClELs6SpeIMUP/L6zqtmLueCM48MqWCk
31i5TtutKE/OTnp4Ha6GRQTtsPOu8nyOS+VYBMONmVe4pGtB29AmHFReDmPoUlG0R+HzrexixPQO
PUQGoWQtkrgrlQs0lrCCwVL3Xm9d79+BHuHmWvJBi+oI8Lna1ye88RFV1i2hBzTumqwlnz5rlHsm
xiabYc0+oNiNzm/K3AjCXaGMQRgaexSsyy7HFwGOWd+iVBvKJIxtEPlkQ+DDSSeDr03bLUuOmBCA
I6rajKL74G69XWL5j6vhifE67cOkYh83up6ft99ebCvyYN76duWLfF0jbz0Psw7k5ZqpFdGtN4CF
8rbcCKpv7DEGtsyu8UnhoRmVv995BWF1dt5GKyugTyzka1R1leHtXr+KWS31jZ+YWPqhIoZ+6m2y
V5cXcq9eEaIQM8hg+xaMUosozxN411DTLnj0gWJuZzd2c7T1hFfxmVLqgJfw7avr9tLjssQwtKG2
4CYxudp9P+5gp/nDrasAA92K4cNOR/jMK+WQ7cHEyGYBqex7yk4ygZCNoSzj8hpUqojeVL0jU5vV
ByahgPjJ7uz/BLooeb0CUUTKWP73LweLaPo5lJ8Lui6qE59pdaEwNZB8Gqajb+S8SX1BZ6wd0II8
W/lRfsRb3buH4ER4DmLCSl60h3pZCMCyIIWsODNE1F1SGXWZq+TFZPIW/n4xjiQ/k/DpX31/IJvX
KYYY9sh0ub+6bnJr/aTXYrpQa6met/eRDAHsTqF4hAoUm035kbw8iQv+7wUQY73xSuMyuAoPtIzQ
zVF0SD3Ev51ol0jeVLGueCEPh0OkuLRPudv4cGyYEufE6Fo2lor0RO+yBLuoJQLQ7GsmIHn6JncZ
yVpw3wv5ogRBB9urb32LSWTbFVcwTeWF0/kjhsxfgj1LwsDp8pZEMEWIVjLrYMKrPrQv4RVMSia+
nkbG3iZHYkXjfgTe7x8kkVbGrHpdaoHcofMiw1nCW0VDwivoEiTxojhAgnxxObTWjq9xGv1xX4kN
tj/6DBgO9ZMB8EPbeMZcyXhJYdW6t/xQos/4LSESZS9kkYh8CHLN8FvixpRFAjxWLrM45iXs/qbC
XmUgEHrPXv2WX51lvbEq6d2nAZ5UUTcxrdirQtpu8sNo64gbt9VmVX+q1eWkTrKKDlfkN32KcDdA
9sOmdr9zJaBAzA0IEQQc6e/nUd0pmRLlIyIgZ7A1ArPPwAu1nVtzfOgHys+jrRhjbDMLaQWJwpEz
WDuqNDiK748cwVgEmVr+wbq9euBAoO22PkCOt2d1MHn08sSRV3HvpQHvETGcI5py9mPdUNgasKuE
jhHeDye40DDQ6Hh1MhYEQnbMsqKLpqgHEdESGkozGRWNVukkSQi5QhVzWwWrrU6iIuXPOM4BAZEF
Y1qh8lwLTEB0j0g3+N43qUHryuFlIlFOn9FTzRzBe/YjwpMPJvsoGRqx0sK1Gew5F8tpUQclem3I
8NF1Kl6ZVmQxaZnSMfe1gfPRsPTvqrcMSW11Z4UCK9QwrV1pWJywRdPSvmK47deh6iVhHOgzzjxK
gy6S6V0cWi5TIXPxFdjCA85ic49Yh9y5EmkDMKUQKJxAdjUzQYs4oILL/QnD8lQNgF9CFKYXRbpa
Ndal1s8MzvE7xQJ16VXcBJad5Uk+V/XB8xr+3LxehQHBjuGz/988oWJzv603YWdFFElA6MG8fNt1
m09z/uGR2XQMSq48YjZGLFl65+D8IV/LVVC1UiGK9zCe9jdYDaWpAbTeCthto96coZEWF1eNWP0G
9Lkbg5mQC5An2wZrVFzmWiVFlcVCjkVI6uEXxMIs7uapLIfBzqx1vOrSAnU1XGhNR2aq5aX2Sli+
lsfm8sfuKcVD9wYFtBuMypDek5fIXa9Y+Zt4pUjHu9zxRT0jnPsRbEClYam0tCy2FRjaNQTWLXhp
bTPNpYeIhd7ZDuVyr+ZOJ9MRGr9CCWBOJL58MVjApNqxL5odevMPnOUO9EU4xkQrT72b8wCC+O9s
Zj/RChQEk4M5Ccwq6PW0duL1Hv2XXoQ/dxUgQjSRjJbmfsnEHhRhKh1HNulUbRw3+QA7VCkyQqJ1
ZUKKwQrsm1QE2Gxgyeov/TsF6/sSpOOWWuh1K/P2NY4d9FHqna4t0tlWbKXoaKLFikkDDv7tMHIM
QlGHK3R69CN4CaqOpKUZ3+cxfN6XNwWRU5DXupC7VAgv6f1dq74SLDtsd8DDU1f1Fi38AfOzUjz2
2+Zeqeb3hvVbZ4rmuQl58ijFz/Oo6ws5DLiFm84r/lVwWC0ciEV3R5KILb6/kIU4wSQsDobA/VKE
Tg7uZHiMdocfLr2Oe5GuFGueN+CjNhk9xKHQyYg5undjawlJ1CK2m/ny0yii/PRLoxgp02S7S0nd
VuoHjkF3kSbq5NySPyuTLz6bnbXQWYPZ9ZGvke22nA9oYT93Z7OvRpDgfHAp5tVPBNSHs94IWNBO
b5JY9EC+HiROuzV1i3p+2YlvdDg9NiAc8hgFHGO/Rt1F17m5BZ6JxoGR9OO79coPO4AllvsJssOO
xlNxlQIc2YcZW4nkmy3bb3Y7DGALaKdSRWme+ycXdO3Lv+l7OSbVHAvACAp+n8xNt8Q30Bb9WQhH
AoCaYyNGX98AnN+3gyzOMrTyY3J2BaVgeZi13/e1n4oHlZFeG7fZGietTEHtaoJSWcVN6S+qb2V/
Ve55898POqa3wWPE11Zin5fs52gcM+EYBH36dBk7Xb6ZAs6v1LmcXcpE5sbPNtTaqdnw2UlMrWpg
GzeOrPRZ5TZyt0/2f0y4GCiq4k2CTNzWH3aUwT4+wuNTQc/xdLvcH69cOixLP/PdsQTXI1lYectk
SA9J6QHslXMI7/12wYQBVEWSdEaSo5IN7k4GU2JI68VXX9FBkKtMBm1N0yDO7ynON3NPhxQVreDB
4FW0NVJL5ue7ksoDwPyl77Vqq6XMqncjdSZgV6C/J+JuIrR/7cMDjdzDzcYA3MzR7aLiMa9MyjQ0
QgmFt/PK0Vwu25vifFMKJ1+frRWPaax05RdP/M/jI6S7Pt5ICJucHl4ty/UrfZFrf5YL5sL6ankd
jSIn7hNpo08gGOAVd4w/pJpYVRruh9ueWq5frE11lk0MEGoxEBFqULOHXtF+iOaHsdiB1jNozcvm
RXhmkLVXNl5nFYkBSsVhFCvDfAcHK6zjCHuPbMuMORgMWTDeGNgqXC+rpiaLo1CEeA5Lau8szKhC
4ZBTaUej4VAolJgnEr5lYjerF14HnfwGrQ+hyU1izkL+BAcbS/ZSFg6da6IzYIhXVuQIIDX6Dmuy
XRGP2owygFevuEhSbhYZN1VnB/sBAFw2XNCQ8AMmAO/zK7zkBnDqxM8ogFlgYI/CBBGQatnofosA
4yNZf3YCe1P/iXgYLH97ZQdkJMUFHAhDzcau0CUJ+p+2wFlwERS3uPMhbzMd4Tb7QHu2UVDtRg5f
Y101heS761Fw4nByCkfDm6bFwUzci43GPtmYI9Qgh3BD0Tt5LidRNZYlSww/KtAVKDxmzCcZTyX7
0QYqnHrTO7mHyBianTDevkNkKcctarVy1gcq7TOOXFuwbd5rSpqU70PpHQV1xqWn0X4oelOxpH4/
FYUZ59sFq9M3l8J8DvZiAxDRfGzDEui2hfHrIEVUr9rP0fEUM8oabCdGLeRyybpBcHI7Umf2ny0Q
wxLpQC5WgCu5Nn6bDC1YQp4q8o5fB+yLjPs9RXV7wvDLF3ee9R6HyJuFpK2H3rOY1kKCX2A2ru0y
DTvkoONKSBkMeR9XT0ZOjSttl+8SQzjX6qqhxoHeLD+eDC2mILPNefag/31KSAppyXJCT+oLjLeO
FdyNKGau5tX1Ye82xNjEJrgOcOT9FaFL4VdiWoTDZuGbeLQEDMhqiq5XOXjaQh74ff9v2R3xbxCI
9N+HsLp2km3inzFiIEJYlAPIHwdpfoF0I7CMZyhzuY2KiE0L8mjcpW3A/yrNwNhLfFbcXiuLSXzP
jS4FFGhsL3OmI3NIFt6bKpHHS8zYLacZA71mfji74pTvzpkNToJlvw5Y/KlahSEPok/Nd5zqj/BM
9JtenbM5vDXfe+FB/5wwOTeImYYBQO4c4wUpQdJ8X81+ZUj/+GZtizqXEtvk3vzznjmYgU5tgn4c
RbdAydKr716TjSkN72ythgLppQ+fUFZERXdNpm3Qo0wI6gIj0gjT6C7aA/OpGZ5Ie69xv9yluR3C
GTc5mCBjYyosvExZvSUZrMbPZW5NPb0GWRwQ9dpWMh729ksbm75CcajlskwGMj68slZhU95sP4q4
fsQBSjFhMOoP95AyLZGZBzjCFjLeeEVEZL0Em1LNJy56otwOZFsE5GtykgDPgyQTM2dUX618IfxW
c331fwCe2ZWTzQ+7P7hw9bzMnKEK8CLdDMIBa55XLHX1ytYkggt3m5y9o0XLzQJ9BTTMOIFtDhcP
2OG5eYPFG8W1vLHMeA+Tq0sVw9D3/dY6k8WlCGXyBNFACF2Us0TGY5taNBBegu9ru23SswEvVtyU
XeJhm1uovugRdUScWVFLI+XTHTQ+mNfiBs/qrKBGH6X5OYxThZJCx0g5DW5HsY1dh+0o07h8Ztv5
JO/PKcSvV5EoIEKhnzYJsMyzNcA+x+qA2TfmnVHaSySVPUYhVg9mLjZ2wFZvSEJWRi6pVwK7530d
s1OHWccWT+l+zI3SHgcLOgOOvXW4xR7H1fyHRgf7rUiHxu6DES7DoaK6y8cGM9AZh1YqFbkLW4Dg
NHzlulKYOVovYkHxrGz/rA9kkcQDfEQqfrgTXZBUsOfTHYDjffbdByoS2w0MCBsGKhy4zMWRMXhE
vf3zURQLh+L3sZujW1FE/YcP5EbO4YvIkogSQQKbGo+HEo4tGwVLAI9+Vfq8alble05mtwH33ukJ
LsXFb1ZrRxPCVh5LQ2zvsNelj4CTPVkyxXT6Vp2SvOtjLCYfx+viw+OO8bkkrMOAlyEmt8Pd8ck7
03TmSMxZSrK3j6aegWeD5B5ZezCy3maJyUMILJ+hPzQTBiMUYaztE+XQv5ONFHj5jhv32Fg0URFF
HX3gDA4qc/E8cYChgipuncc389ffG71i/A18iydmj0MI8DKGwEnlKXHSdYyewMOuy8z7kotR1CgO
NiNVwjNBtUpyn7n+XnlZSuQReaQKGbA2d9Sv80PqvNzzEBP/XHINEsGjfUomtn3vjxbMvUHjYWsY
iwhdUDB4B48j0dxuExNW5lwSAHiQu6aQyrX3m0SZRKGOISA0rLo+UQxTtKGQWfnteAxSwx5Yexs6
pZXNqGOIFrgHC0mRz5aZPtbIlSKT4XKvLdATUkiomdv25toZvadDRnTn3CdydQ5puy0ibQ/o7v4p
ijz1n6Znqwjxzajl090WMNcaEI8ZderwqMOU+Q7ARGXVJ4gGty/lIxXioYZ1kNlOEoHzRgqDpSb+
EqfR1MKB1MbsBeaNcMyhKFruDtaHvclKhD1vqhcYmg3AnIjJYVbGcL9XeCQtoHK+M8TxDz5nm/KP
5aWo9GbAiEsup8MT/4jHYHUWSh9Q81ZEqrsM8BTWFYz09eAdA9Mpg4Y8fnsHCJuCFTmxoQyMIU8z
PblhNs3/rq+cMXS2Hxf1Xi5I5PjrKWsW/p/MzXrqXJBunnlhL3gwrM8oEWjgCyGGjPBaAJNCKSSb
RyJvuV7p9POdMWhhLt4eZ7beSGZ+2x1in+qWHXLwAHnzCWrSLpwtRMGQ+kjmYalH30um11M+o6xQ
BASjILIjzb+jZh+A57qY9qBH/gxJUJ7YAtO2O4LT3t3YFtxRFhA9mFYsD+lxfJd+p2nhKZDC0JxR
fHXrrXBpCBVCBELXGayhOukxPVaG0wozyDX2hlTl9Q81GFP9xr1vbbTL+xfQ9VDrPAO4kA36UtU2
/iJavS/FzKUF3lMG+h+X8VBmng//NZYZWwv2gbgR2/Q9Rdilu/7MnWvCPVn1NEIx4hsqMUKBtxSM
yHsg3ee4PL2qetMhLA0IWWlW9+OeLAGPdGVGwX9NtiS0LvXdtHAm5PG6LmTagAvI8xH7eO3w04SG
h0q+ujtyfAqqaczPHWrv4SGvIJElxnQlxiWFHGZKxKJftrbYON+IDbL4i/X2rFOB7kbfirVon4J4
M0BnEvkfWwAXN5L+AUxm4nayG7qQVP7C370FKDjuz3GRE7YhYcG5YOAA2xYG4Z82UMTG2fsfupwC
3ZiLZklERckeJALjmt4F/ew63D8m042h1PkOVv+NcC78GGzvQ0nZlwGjQd5hdTprGG9/QnLZ10Lc
xgb35zq5eDtiUULasGkG/uxFGn4DHpLXiwN7vUVvKvxgrv9/vT2/bAO7KIUM/PLQcrRRknfbQ2Pr
Gf5xaa5pn9DR4NRW0Dwkd2fWqnEAb08JTti8mGLAKG04wjJsbiHTfYuTCClw5unyTVM3aCeaCFlT
m8pvQrz9VtcyhWkP0F9EhGZ/6f6q3RlYe1oGueVvnhk4NKoDyVL6r9AmgGuErlYxCVFux8uT+3ml
Do4K5VWdJiVJtoNd+VUStCcJO7rzcJF8EpSgYoqlIQq2pmuh2PVFo2U0WrVHv2mdOz9ZeebNYo20
QEpWbTGUx+rKdhes83J9XIFkhXq6gzoXg5KgCcltuDGy62wCKM+dmiGHwMGvF8jPPNad/rlj0kO2
xUHgeTGIkfPmkaJKCpDcM5J77AsdOnU3Gx8MdyKXPmyZ2Fnb9qex5IFcRn9rULpWLzV1KWLZFYHq
PPMDWeL9xAM8IwEU5gxN7YjVXkHfDtD2AVHnRQ2FJbP6Vya99iqf/ryCpxbS82cSBftxkuX5w+96
mB5/2q9DgXEbrCgSVazBsmPss8e6tg7neUrowZqEf3pNyLLe8Wr7O3X3hPzkqIqMA8PK4iKO19kl
wmGBwnb5obiHpNN+YlI7KD004K+mi8RN8M8c759BPRlwDDbFvgzTG4S1j4gQY5RuTGnpReq49CFW
+d3483bRdNcAb0b81ewRqi/bmPeg1+UIGLbIHouNwYx9o38b9aK/DKs+IyoGrFzKziDhzHt6wu5b
pZJHs7H22+87zqoyH55CfEVBJz54gfCGX00njRg4F4ccWcaCsnmDTkDYBORQeFkdTrolGj0VIPOj
/6OjTTvg+8liddscZ+A3kSKFPRyNDbmv7+/npT/K79f+CSWYqTyzyVGscwf3OPHsi786i5jxc1cr
1zJhFdTHjqHsE9hSoUfm0v9ztYcxSZJljvCNa0mIN72ks1D2m62F1Z8elAAhjqxyn1L/bDp4zrAO
tUgCAFLaLSeOmmd1bvkcZwAQmBA6x7+cw3MF4Ls0kYAvYIXgJ2YqSmIxjSarwlYRzAidoFYM9dHC
sn+lH1ixh9B2Zrt7QoOXTarJJjdQXsNHiMPodJWs2IIvMF09I+XAKN4mHPxOpXzojS4zzaU+CDZh
IVa061zE3qypCm2pQAHrul9Zy6VwUcFKSI2AnPdoGiqyIXE5CvM9gXQjqIGvwpy3hMhbFhhVQxMG
xyMGetLicVTOx9gwFdGAbokxfHhkviQFYa+cB4XD8QNUEVjKoV/iKbfw781lLdKtAz22EXEsODhJ
PDn4QEshOykJvFgVfcq9+VW3AByZQ5wQCpbBuBP451dW0UM1HBDZjB0K2MfcVlTUk4rbS5zbtKja
Kh2NQtvXq5v47g9CY1bplQYgmFTAFubtdRXb13uYJsVqFpdgOkehG+g9GZ63eylzHTKkyvRHh8py
xyr9wawPc9h4bOQBwzqm4YBWq/p5vQuGN3Gw3Zyz5/dixOvcaIUyc9hRASYvWCczDhozLSRYmXBw
ppUJEAXnFbXPxKrEbaKb4N6ZqDdxEDctz0R7LQ1aHYi4aQDmajzgp9GQCPU1OZ/H9xDxODmoiDxY
Z2VQVKX052Sa+8no4Jgxp/FcqpqajhErb4r3bkvXOv39yQ3WLrls35YfveFjQ0nWeezBi64QjaoV
G8yyn/R5HZbp7C9EOXPPb+Z6OSYPau2ytL5Piih0+qhBphh0aN5L9MOkTLalfnylyJwEGN7VNiph
KcoFcKjgwgDsWrEfhN548FSTxw6azBZg9CBWtgvIcU1iJxDwfB5kj/m9jA8h2wS9VqJ4eiYWJv4E
qzZPRjFj/zerMpbWcz0HCPNkRrDvEQoyXJmJBLi9VKPK18DFUZgs5lBmUXTA8r7c3lbAhblLFxY9
CVzH6iEGQ2DdgBMvIzXa+aLoK7itBfKuEaXayKk3em9dikZHuGMPCwf+eQj7taQY7rUcPWvxt5mm
tPB4keGY9WQBM9UFHTlWhcD+5EVsfGxumKq6+2VksOIyy1uXCJBrmE+0/kDEFDvsc06VSMRixZEX
mKLFM1H+R4mJKBwmUqXz3uvKxEJjjDfH9gqWMo/ZNyMPp5qd75d6dUpQOjxGF7fXvNIUtLkA5CLk
tGS0yAiux4X3rXL8REX5RV8U6IQZtPl1Ag8AwPiFOg5ddJ67N/BeXL4qRTj036HrjKggyloZj8p1
tGE6hh1zudbBXFq/imzhzwfY6+2yfjxTHpjFJYNfxNU0WUy32UVXiYzHyrL8UhPK1AjPm6pD2NjI
rwRbBWVDZlc/p5uiKtgmnfHjoIxRoG3oyBK3fckvlMiSYxbm2/XCMJPBM++STXXLCrrw4mkBltjL
W+y37n0KjXVRukHoi+P+qXruraGw0JAbIs/ZDjkKjlWaZ1bMOmGfkuaLzqZSbYSD3Tdsn9R+erTy
Ro1Kkcn5lJrxNuXtM+J+gGsXQKXKn9Ybl4i/WejDP8COBICUOvCxcm3cNxchIDYeAHsppMxtkMc+
STfIWmhWq4PfqAmHPXma0H2v/gdf+U2XdZVqcRYnpfErdmVdKP1VBCLsdoJZgD3IJfJH8J66c9Sd
WRUeazrDmSZMowjHVZ7TT6BG5sk8GDdKX9k7J/p9PnC6AYpbtctA76BQ4mnwokelOZTE2TpOT38A
1ygRpP39fl3Xx55lfyaGO+VyWUHpBJaTobyz/J0ElCWTkyPflWxvpTqmIuE6OglpSTVMjfzjijCT
NzF11Oy9BizERojB6L1siUc1SPyfb8mEoxszGWjiECMpwcYDqAKsi7nVSomG1ZhzjC55HOPmVeUf
yS4a5MS0ZuuNij6hOx51qwxJ3RJ3bd0qr0+Z/ICN3WL9vH0YxTrXh0U6mPQbBbAzl3IhTHbNV92v
N1lfTj6WB0CzNu0kUbld855zbmpq/d61kFka9wj1+kOaPXVEXh96OoOxbjb4oTkpnQeLG5aai1oz
adCspVld3WQM6yx6pWBwYJ9b3eJNRER64sGg3ZgoJUTRyBKibHlnD6bYReaDEGFImNx7E7I7Msqf
oPfz79pK53B7O2L6uk7Unu0yFUylPFZ1iHVwYWflBFrXIBrGu+QSAu7cS2deLCZU4i40K+Ky/eXo
ni68iXXqJBurxxqJBLez3Dl+ibTaMGai7fwYVfNfyNVGRl+jT2i+qeaDZqFVo8XQLvENdy2U8brD
GyGiHCsPBxv5y04tl1/cNlGEFW8IV9nUTg5zy5GkzyM7nzFndva/gNVBuEDjXiWZLjE7vwvAt8Bz
+vmaOBU9+0MJNHbL72q1bUDhQdDFDnbEuN6xpBuxZRVBXpDcCTzc1fI43fAotcdGUuY3MaulD3m3
zR+JsUfM+2aC3rfQ4g7D5TR/bDYcrk81qfXlgEMB7p1pJHW3iGx1jsBP3ZwaffGluvMVg+z1egvR
2bRtUDcuTfEpCnAP3JSzU+ACKXF+2axDBbq1EWV4b63O9j1K8TyhJdSf+7lIdrPjpw1GOwwEMMM6
jc2Or1mz7snMSjaREUK23Dr5JS9bD65eqZyZY1Xo6HCo8ZpYaEZhjLW8xdSjudjtIQgGsDgGlfUo
TgAicl9Vbsn4AJUng1+kIOqtf2iERDbVe953zwsJgM/Uet0RdBTpOhJZMcbygGUBvordMhUq0N/M
v3fFnuRQHHTza0Eeo3K6vVdXe2g3wq9MRK2vug6hO4QAcugDKiZ9n0VORBCPeUT+ejM2/3CFtfuV
Yxo9rxMfs8o9aClw3whOy/Z84/f3Tc/YA1HfHGLkMYuat27wLB7auaOq8LFy4NiPsA4G0qm73TL2
19sEC31ltWsZT9eV6oRDriEd69xwQNXgGSqx5GSDhrBG3VdFLSUwSCo4/rCN//mYG3gJCzeb7TQ2
aUdmuNXLOGzsPB1TAv3mRrgKEWjOCgLa97/JXZRv+4+rqWHL4EuAkChrOnFMoNNQww/+q7o08tkl
mJSCPDzCXfSigYS1mH2DLsQ/pv1XtesxRJj6ooF+jCufjDkKV4sBFynakpprVB7soRIDhxCpZ6lj
WjR3TSkMT0ty2eaqWZJXyFNTLivbaQQ/vu1Nz+4HCR+ELvzvrAztqQw6zXd1DIModpdLTCxIpOOb
UkkR8xFMb3pV0s+ltbYBlPbGU8KolbVqCIy+XVre9TLWh51GRcgaEurWsdztJGi7XL/C21GRytGp
dQRKWAnPQ5TcKCwdPkSM4zm9+k1kQRcNA3TKXTc4vngHAx7M+Vp8idlKgOtUEZsuixNuYTsg6cQ3
0zr0WYrjh9lPmgcH6nNBdCSB1LkH6Ovqp0F+Jrp72WgBlpqQ9KnlNAap165XjP3jV/uJbllL8CCy
lyM8GdmY2fUb/VVWyuPmuiC5rT0VKFHeSmqoDB98/iB4eb08kcsJG4km/tCkiO6EuxUzLLhtw4Zu
4R2IrFOGtAUBcWzdJX4MYSJXg0txyKm4gNRfwaYaP58Z/X6zlbd4anhIdEvHoqmkqF13VLsRuZia
kBuIq3YcQ/qvcLa8Dn9bQcOfF7uQb/Vrm8pmP6lg/ZfclxxUpnHwzv1rvgDiZWUVszsXmje/Xf4i
RtzYXfgW56cmZK+K3BEquAFwCDb9lBRw6QiUIimEI0OYrMPydGvto5TnNdE0HnZOkCTav+kzGnkR
Vk1BZsQu+j2maE6MzAOvRVK1VZbt7EqZ3atfLEPgIC1/X+CPTOo0qNpEnGVsL/Oo6Zd7uN3KhrIW
Tv6fh8VPzCVJjvqljjENE4WFv1hW0Enpnq/XGEcUY0sPFmNnwXhEVCIBsqSZ10N/ZRQVq1COykBg
+dvix71/bk9nAihAo84vlYDqJA08E9bR5ePQ80mD1rZW2A56x06a2IEURyHTEWZ+bTD7dfFgcOlJ
w9TsiIV/2kIHDwPRFsqztzA9Kcxp+ggwv44eWx+KYfDLkbeKJrjINp3N2h8Oziek3KiIBKZR41YE
wbC3XzV4Ku3/gPduJMeF2GLnydUmYcmkjHoFsisUHG4lmT4fTSdn5byHo4RrmYBhIATVis+EBt0M
bJDhucn0Oah5JyIW9PjfD3fduxJhnA+6pnsWoHbFhsVu8sv13fQfPY67PQHuvMBU658wO7fqmmzN
E5jT+2MhSdnjU1a/BdRSxcYBIdmJiKpu+ZHEV9lGRU1LUgf1psTdcwu3BefKEw/1PnbNe0OuBu5H
U9+dXLvwWnfRB2Wh93qQKpvlM6NqsnXbb3dNBwrb2PxJQlHQaDEOBla0ENnNfP/+81mm3iCd8qew
M/tjAzmk+spY41vvm0r0UREnBPrRklGbQHSYKVTA091r0jt4TujW0c2CKv2NvsGq5Mz3TK22V/YY
WOtFM9POGQht+mB7PiJIjjrLKrMBggQj8Yxl9mW0xm2h8cZtIg/qPWQP5gP6lLY8/3HXXS1splAZ
8NVu3IUKdc07uEGUzXyctFyz9SWuWiA8Q6ElAAQs/5xp3VlV1+U1Itmhs+8B4DkUtsdrWd1056Ua
hYKWlS5dwa8H6GwMe/gWopCMQJnlTtuMYQ2d559lK6rQslVFwSDvLDp1BbL9/QBIi1+BkdjhUYv/
AWEIsLr59oHEOrNc5jWz2ErlNLHrmW9jFWXZZqUjbDl8x3NcgcbR4FqHmSY4HROviI6YRh1C6HFw
buc9OtHjOTLAHv/eRQg+e7tZJKnfED83BF2RnNAaSfI4ywxJW6pNM8rMHbaYi2OoM8F4mHsXHSG3
4X0H9GhRrPD9T76/ihjxjNZ3Ye2tzOB0JnIvEUzgAnoOdBnEAOskZ8HUvN0UL8K1FNx0EQPiWLfK
jIi+RGW8fuTDvWYNmV0GlLerT+6sePTy8YIpKXhGCeG0UGyf+Fl8AUZzUKrROZ5bg0w37UVfuCl6
xgkgB/RfHnFCSESnIFd9YJ4Dn1C9/3hWwhdwcX/Qpy6hrZfu1Os+0xHRH0bJWg4RLe7Qqpws3HAE
HamOXvQ/sZdPRptheM7z5cxX/XY7S1MdzRCTMjhjEociP6uRsbdlB3j6TwFC76FYg8MAwlFdrhtu
uZlq62AaQCkujaNyIH2JXX0EedAxRaezfUJcyr6PCxC32MpTV6jnTSbIpUFMFYz+t/ME6MA6G5OQ
E3Hn9/zpm4wCRydj2U1sKMJAk9vjks2EwRZ6nf55Go6WjbOnfjKGm5siZZPu4SGEFUiDiFaeWNXv
+yeZin5wgrYjcPj96QMXTtYfS8S8oGvaTDa0b9kV+/VOsDj/MjR7nVuL0dWk8mOakugAq6QJk17B
abwy11JrB+7ifAr5bUt2jg5AGNKj1J9pmkPz34za2A85xOIleuu5nI65q/Ykbwcdx3Fx0fQZG3dp
bqAbThh/m0AYbhISobOp6jQJUkkcMq5V/yswww7dptSWDiSIt6LQSD5D0uzzKOXs976h/ALhwVhi
og0AzwIT6wEnofmrESHqLhvR7Eg/PUTS19u8kMoOsnVO6ybhcSkEGVGcKDh9b+hjT4twz6IZNVeF
ujSUqDhkPo5pW+w82jRY22eOXUUzHEjPwQk3ylIJ9OXmQxxVW69ArcD9obj3XafJdXmiHSMNvXLm
sb13GL2XGk0fvIbG4DxmxGXovu+4Qw+5NSv/Xp5ei0A7LkamESpXEnrbNHuwgc9pRXFhhluyyfxT
vbbZ3L4GnSGXKvG4od3HJO3ipKFoyPFm126PCfpr74s49FbrZ9Z292BIlDR6eLz+LCYCZR/W0XY6
CQRvF1DqL2METqugJzm0uw9S7e3PuOjl2EJ/8JphbSnZW8RTl1qCEv3oI74GP32OF5lr02SFGjXp
eDm5nwknyrfi+kR8Vh1j8H3Fvc1Hbbw8+2h/gnTmjcdLj2YuGe/tipuZ/0qUBG7QDBqg34JCycb0
43mlapjTr4Pen7Rhm5f583w+xP3UCqkVh659KRQ7YvodUo6+No2ItRT8pf1IKaYO1Rot/NOl8F9S
E6RIdqSLVm8UupBW/JgXckwA6j+KQEh61I4fspOHeWNe7lBm8AeU1AQLPa5CpEnrPH3/5dckVurD
962yxiznqhUjbZk4ohwkSCkODauZDTOB8FYv3tButxcb7YxYTCgsS7Kh++GvsmJ/PkaQywhh+afv
eT1y+lrXvJLkAeE5YmS0v00vHzoGXZBfUGH4KM5FWmY1rb9WiLk5KoYj1FfiTLxLuFx+vGwCAyoI
3biXzKg+SfLQWD1W/iiKGmTxY5AniQz7SuabNIzcP61M5LE2gWecvpwUUthqcdgIbUelh/mLtbIt
HJiWwEMp6xX9Ufg1XHPfJC8G9jxGS+pb4YjxnLmccg467PZwc+XK7pM61OeX2z9fbVDEDowR5vSq
uBEe+2UPRIGakF8v+qFvOpgPkEp0CmJDuIOTOY9EF19xRJmDO1Uf1o/HXcajg//vOc0HrJIOtJJn
Y1U0eyNS7xlKC0SpW27I02F49actO657fAUrQmP7U75K92VJg9EqFXxTZM3fs3M/dHWjfAFE5Ek2
7d5NVXk0VWT1npupMEcrp3Pl0phiZouyG8uvXjG1U3UmJ+uS0huVDnRD806B4M4Vkyd2HaVEkbCH
QfWsf3CrcOTPXYk4hTZ4WMb5acpVMnAOBa2UklTnLkTaDWfSw6Ihajl8xiIH6Qum8SdQd0/6bcbQ
bzG0Vh/tuZOfX78e7QZNY+rqcX0X4/PuA8y6kbVS/TCNXqyxlExfgia+v8KYEcCynPix9tZEG/WW
mnhl8ynjMAaviayaPxgrvmfYCDmzBkiSC1Cls/5cO+sNJeY82qbtjbP0SJ0ljhmV7ZEGXqRTNT1d
wisVDw/4mIeRRYvxdt1obWjmfkrfig6gRNEiqlwT2PT1lBZMncOkwTF6DuLVqOgusr8sP7bxoKDo
aeoY/mtZg4mbexq31DaaoXpAoiURCo/KW2GGLVF2+92YwLzzwvisK2M1gfRMOylB2ke2q2cIQah2
Teg1edFt8SWb6tudp7Wl7scQwfoCR9RTJXVNxQsjI6MUWh+kC8+yPUO72AZR5Vj3zf0C+KoinAid
OpBjMAEYkzmoAp4TMhanWvpJQwo2oGB/SU++OEqffVSCcGfODhwHAhDEkihPq9jvc+Lxfb739f1X
OTmwhbUwSSA+M0bWqS3TTmoce2eoLZ2zir9I04tOUO2ZZZppw6BuSo88QXCVh2mqr6k9tdbxEYUC
FcxxpmGYrvYzZ8+IjXFWCm1bzr9JWsLo2i6P5ZTWr4jL6dJs/JI3fSRKZlHbujOnsqYCMmDZlPLq
mWnYMNWK6whForLciSsvAeKW194tDyxWuNrIVBbibp+nVG67hXIzYisJnvaTthI5d9GAxoS0dzQo
HAWtGj8/0Ego/j0cJ+tk9YLqu+I+adEzi4L+FHflwt93xdDajOAt7gvqQwMr3fGa71YfCELVRcM0
W4gyjYFq5KFSK/gscvcMmKKG7N8JEYX19tV2UiPSmFG10IZAfjaWoTugq6cy5Hmlcwcg/x+9y5PI
fvxV+zGLtSwXTqI1UKrvetiqWoQInevMz3G+/pb7UumDecKVd9TwCHh+YfjbwEy0c/X+TKRpQTdd
v9W2TUA3kNx+mZ8G7fAy5/BZFouPsrh3O2EIfnTsYSQvZcr08UA2y2izdQ8+tJov2QxQnGQFPp2T
8u+q6nz3ugEaZDo2VxRQ3zre9py09l2h875caxwZoyzSKffRpTyvf9IZiUGEv3hngk2C910FK5FP
F8XUKPHiTPxCF5IGNYW99MpmymaeH9KzxR2i0ehkGPJOlJVgNCb0lev5WHQ21Knu7LVmGwLLJm/G
am5JKluVziG4n7hv2az6FLcLTHC0XVT7dicrJq3nrtWAmsSM48hD1OjEu6ALZcF66JKNWXaEY5v8
hr81ylFwKMwAlR7Brcrm8T7AGXHXeh28AZ7TD8dB9+C3SLz5dFN4H/LJP11KXHSCAIebIX+8cOvr
70P2VxSp64kz5H5SxMIYkHemqA6Qhr4f+eg8xDAj47Kb2h00KHUi55LDF6lCr7SFeOB/Kmfkm3U5
ewCONgobj1LCFdmTs2whqpsGqGDsxqb98CaXYUoKq875piDDaHlFr9LXYjV5HYQGLZo2INdR21Yb
dVjrDTydws0gg0Iu3IOTR1/4Iyhpzi7iSQBUkReazDrhNhuOHZHI8xOSGEoZ38QwTHNRJQn5zf7a
/cHeYLxaXriklIXWaZnaVMId1ak9UL63JL3I64S8uSeqW/yHrC1Jkbigh2O5NHCu1Bhoblyn7xUx
zmQ9zq7LrvPlGVg/pmxXyger/ZRNSNwbsQHz/UPfBR7ILsVxfcGGEuvHTfzhVUNUNY8xMLqKafiD
hqiJetuI3HkWws8lNnL9lzoLB1wqcLlXbqQsJsg6UEod+P0FAAt169uBlGaFWn30L0sau2WaWAob
5AqjYy+iQmfEydxmqy9+OUmvw59GkTfhfnxza3ia41AjE+v8v+MaWyUAlrRl2J+v7bDCZeFHq1JP
k109i8/ngtglXopkSaaqimMOqCcR+gfX2UBMkGk5SyF9CjhXZvEWLdLBk74Es5HDoKSnYAxmqs6/
S8M71H/G0MEZzHjLnJrrq06wX+ENosiaLChnSTP2ZexyJweuBXc7uBGFnG3u8QYySzQCdj9g0X1C
JI0EF6zfihliJPeUYyunxnvbLcVe2eQrKmXKPM2aYOaCLr9ouaRaf/gvAELqYMUBnnFqVLbynW3E
oHXuEVb/lF7vq/MOs8kZ/xtKaDRZ3go5qefCxc/pSxSVv4f1PfkOCRHRf5lBxfaGdGIjnMbwuQ2D
swN5meUGpmw0HUsZkjCAY/wyAJXVR5jkRVPGJjIBjmvOyk8u2OstCEeNRoWOYR80uCCJ8MyDed84
u7M+8C7Yv4ARmlkX76cxQltWBMNLMILAF3iDzIoyp8MW/d4CtIvZnUs2y8mA38HZpzQn5ecUgyib
iYGEY5OvaYPJFzq+SJQWH/odwZeneWMnKnsBL9MM6Xddbm8sxajZaLrAUUfF0eyJjNIGJz4Kzaef
Xz9ScgNJXFHk4fdWdqyz7dCz5zBWSDip+qr4TTHI0WS4jG4yJXxQWG3Cxuvb6c7eqO52w6fFp8yd
PRRHa2druNO+T6MsWxljOh/IldRJkOnbQvKJ1+gZpCU15ujQbF8Ze16SWjiJW+4CQzvPPxSrVx5K
dXz3XhWv/LwFdclZn5Trq6x3KGfCkT6ui/Dmyz6wyXesXayH1wAvwSLixMRy77qLn4TzS7adLzpF
q5ARuf1GeN71YdjqX+fXDQ5qORSfw5E++s1PSdHpqAImqkXODGMiHS7owt75MT3HPU58CgqonxU7
455KBkJidaz2E5iNn+ikskJ6S6BEx0YGHcQdQt99k0pRbEwY8GeFVYo44Agous1PcWcDm+ghrH3t
E3ZQJpe6VEkpjFzm+eWAMfszF03k6u2n2cCkPLZwgEqpLhJauYNH6BOV2f8gaxRYPuOzU64Ui7BT
KgvDdNx+TiCdyYkWaxs8m/O6x1ejrOj7t7vqcpjASeDrkcpl0EFXwY4YXvCs4CQvSztOG3DX/I01
YcJZ5+fjlyh4SnQ0elGI4pPC0zOZl9cO8LAI8F2I+ABpRlfy0zNjwKNA6LIZMLae/PrjJbqFP5GH
WwVWXBtprzVoubpKGStefyEJJF4WY1ssvMUQOM5EO5ncsNVaJNBXsazejWDOrRQj5/7L8x1NrYXp
AY2QeV7ESHCWnqpymAFbMfXnuFvB22p4IJ7MU82OSnAoL+PDD+40jKnE2GIWpg1WCjk+HUSwUAvD
qzBa1WFrlq55zDRtAEXu/zYBKxEqNE9nPUjIpuoac3deH5tWWde6n5es1I37Cqq89wP9GMuUfXG1
TE8BisLpWPM6FBu3WlycLEnXy6U/qRqx0TDilkLOqGemA2Fun54a3N0JxoKdEC8GQ4mLSmsm+WlW
Up3GGtn99ZKORuyeWnI6Mu3qj6LpZktRgC5eHDYOXZUjwyLRKirUqLG/xC0KN+aIHVNFGKmrbsNH
/MccRmNp1L2jpmzNafH38TS/3PQPkgoGLsf9KpKb+P/K4pZS1DLCe2Jn47P1KTR+vwcVMN7TZBvx
XGalc+RmjHMMijBt2qO7wLD1YKcioR0L1s3M8jwdJrE8YwP28arS6OX2yrpZVGGQ2KP/pRU4MVKS
iHSC1ko0vPbthz4PWVxM0MKLVj8Quy7k6a5h48PdXU8caCdTpio1n73l8LqhPm59W5GXHHzvJKno
yXJSIPuLC9QSCghmm8F/LEvT8OrUuprJUX98NRcg+tDl9bkdt1lXGQ0dJSdbAedIdPkUiiM1lU1K
XrSS8es/8lWvdCCx+kQVXqnR5h7Xo3mHakW9hc2o7R9LuBBrb+2fwPOp70vFEouRUVeVAhpYHP42
NgkOKIA0vmcvoNEKcXId85lPNugNe+CYkl4U5kVk0O3a3uYDA9EL3c3SykF8Jc3AEUnGOO+0XuHd
UyEgC0VKeJP1ZLGIP6ks5rxCzinrhdT4jFWQzOGMn6wqMwRV5kVbLrLHMJaU2r1urORKsTORbEnU
HYYS8rlPuLHvjZVbun7FW7qv3GB5Q6vVdj23Ex/SSRdCLhJ4FByX4VWoXzb3WaeAYJim7jfZYf+l
bQX7GFIchPbtMwvyQhOqUsiq3P+KHJga1aj46BYKKyds44qU81xYxlNhob5Rm3v0/7eDE54PAwaX
pJiazO9DDvmzCMyBsg8otMIpWxGQtNSF81IHlQKTwP8ablUwbEffukCURKF+mq99dy/CytbX70e+
2KDhuDOO+mE88vxgAVBWdeEhhk0fkmwrMAGgpbSrLmkNykXRxU79rkPovDUMusvacnILky61RJnw
e4cwSLfw9LTwRXl4uoGneR6g/+OhEGhcm4ytlQmkrfyqvbeRf+fS51GYa7gxxEKGRqdKk407afjz
kqD1L4XVsCVTfWsEAOVbyEmyE+hjqgeomNSjbUnH6HgFuukqvrosaXaKDCA/fQt6hctfHOu7yDPD
q6yctal3VfFq/vxIiG2/4Zv5iqDERcW9rtu9Q5t1fe8jgN1W4SsCZyVUYTxVBUDjN0367nCmkQuE
436LcMXs835MzmBvpNu+NXPzMVyaKlyLITmqB3BO0aGL5Dg6/qVkuD7wylniee9tkzRwfyvIhmB4
KKy7EARVt0TWOsIsCpGa+U9QkDUsNpkCGrk9Kg5uxogLWyGTwdN4Fn8C5oOjaCdetr8RU+JAOh6W
k/shmPkVnX1LhonH1YBnu+krGvZVo9FfPe8xlZDRv0p4JHn8y44LcZPSyq71mNvSmxHA6pRk1iCC
4IhnrnxVP2JqD96qZbedpppxqHR6Hb6R8NOnELZ5IaGIdpIZ0aktgRaPA77IfldDqH9u+Em9GMbN
z7amThCGX6JP8KXVwVXpTIZtpOXnPT4+xuleZKdC1ZSJDtYblDGCyXVzsCZYiYWQRVksMIAECXH4
SKSU6kQt4/mPNM372m9Mo0Z4ZoD7PTJE31sh1yZDloBbl/8NGVotwpzvPnFq0t7wosGf6xqACiGf
bThegPLnE5Uwz9AU+pyhi+8/HaNF8fiGYO4mBmUxpZFWch4WOHMXkZf2QkCW3zrvQJCiNnty2673
YdRlmH9o6CD4I+TLixB+xRRcBa5kK85gC5hr5WBj/rnKkVqya3MUjTHSJTcMx26kLOongxrUN2ih
AwJmWU328OmOL8TaJGaF9h0yMP2W3fIm//UKqtrrGoDnQlMZhKHgV7Jg/LsDyxQ4TZgNg+8LxN0P
optI+Kgghg4w3Yp6xDSsv4z9HYrsBUpzstGh+3GlSyVirG5IBiAPa0J3/mlMjq2+hndUGUPORf3K
gfTpQ2at690UxDrXVQZismuGFhuZ1Jd63jXb+06HVj9CFKI7L7ckzRmajZA5e5b/LJXWAMtMBp+2
1xrOVQlc3YNoq8T1JprGHVUjx+WNloEvClwLV8iIh74lIT1dRxPgfuExt+1ZJTxbFHPjlrcuh/2I
PAdcBGE+W1Q2krpDAji1nHWt8JULGKg/Zl098GgImbgJk2TcaKcZwu3W4Ep8jwZ2QotIEKWeB0uk
n/tcmjdjgLYPZMuFzwLwixo3ZANyEyYvCEDmPAaRQ2euOQ23bNZb5gr2lA5nZ2rNYwq2bU/7R/Yh
Fou+ueBoqfku5IGwW5+2WlMt59aQuCsAt4otD/49Tbo6MXg1KdNC6hS+E4TcnbvCnElmzosvmJLN
ac57+gu0ADBQSMm6c8IYqVT0/Dp4kg1LCnVuU+5V+DteIOkl1TET/cEqYYZKIHOcCOGFeybD3L4R
/r4VSPP/6nzfzYqBBP+Poj+tIgfBdl6SoVRnCegKGUheGFKI0uTxOStOmh4a/5/1ehuOhuCrVHEh
xA8UgSDaBikMLPeTeHPs3KrYgyQJv2lcVVlAi6VK8+lFD8T9TRzHzav0uq4FFby3xvCBUkDCWbPG
TY5Y1iZFeuXapgVQGZykzUerD2IlWlevNBiNVdb8mwxJ90KvnDukGYomFg1mI6v51R15osd0Gqnd
yoHMcIdbJe0tr8sL50UfNlmBYdmy8WqFflWTfWNhAt5B6F9EsbqUJY1pRlbsUx4fJihqMQ4nsxov
hDJWKOiZ0lRycpkiS+JGBYufKrC9xjMD1ikUIK2IjLroWB0mdbEDHtj5oVkKwztKsqjt+1q4KDOE
wvanFpuybbnRRX12y6DPHoPtsWTQ/74IDvWA8k4JdnzYe9xgzI+S1h6tXttvfQA5lHPl8Ol/Ku+H
wt0zqd3RMshufKc0IPJqmQwniJjoD2aNL5fjbrBF7asEDzua9jB/n3Vsi74nHucXfB/cY/BKk/sr
+S/DFH4ztVF/nWyk/ULwz9l5/G14Z2gAlF/E485qneG6TgYcKQDCc9j4QxsbhBAqHY4CxoP1DQCY
KjdX4clbtcyjdNTJCtNeQgrrFTso2p7l7dU2ZtVUgmPaopTviTQjwnlev5vnuO7K3GINlgR8UQA/
AqhWdjWM1pDsZKQAOcIctgvgAk787aIF4GJbffbMz4obTCGaEWq0M2ai1czvxYmStbURl5dS3omR
CfSlVxV41X3JPdBCPi3ZOapWxFbLd2CottTy50weJtJ2QZ3pZAI7oNE+2zBAcq1NZ5Oxt8gzaKLc
dFUIe9c/XqVOf4KmeTAkIoEKge2KHNzloJR3OqOzQnLJVkic0d7S3dbokp9yYgd9t4Pdqt6ZMU1Z
pDM14L7Om/o4Y/JTHKh+VPScdpaMdXRqw8D1E/Q/b2HtwQFCzHrAN+DzxLzgwuxsay7fU6rFj7il
ey4CNAR4iiYPpj2TDtTdfu/0fkm6S4wP/9gt2M9V0Y9pEfVyZ8uvKzpxjaAOX/xbOJAGx2Db5Zmr
6cAbgqpVE62T4PdbugGmmgMziUBcbYLp+8sl7JKC8V6ugf7sOpK6FYStQRCzPx5VZBbgz6Mismem
cksOTpIHh0PNP1ynpUNJHXmxCCluPsyq4pLBJg29LqR0/9471/nooPFeGQ5LyfVYBaEhfr9KKsH+
1o8RQO1BotuYI8LbUuBv7TAExL8l3crKtOajknKLJ5Im+S7Tk1oHNYUL3idE/4qdR5Ni7FPOauM3
ZU0SyT9jCZcIZV3PqNcAwr9MAwcyPxSNDssq9SL4rtjgAmsMnETyHyh8qQOrYMXuCtFNrBmuYHoG
2FgkZ8uLcnsctDWRokSF0dCHe680aX6Ho2JmKPMccV1Iw/64rcvfpIMeAouRoevHmVn5iVt1PubD
FXA37YI4tpnRBn950yCJrBIVjOu4UV3q+Qagb5lEpKAxaPL7wxmmE3WsbgmjfzaUvcY92fl2vT66
si3vx37cvmj6jJRd/Vh9Or9LYxMiZx3FrTFXM4h0hfWGAlgPphqgGrMU8BXkSnYWJGmjhjJNO5ey
v1fiGQfoEA4EXYpJyd1QwItu02i9VVTAxJNQe75byiqmIPCbka31tCRaofbRDIvzZh93p24U7Ko/
+IglFhi3ARRW/Quy93VWJwWdJEiRkOyOI9VbyuJ/JvDVyjGRwdXtPdjtBsRFskRwVRrte8Qsnx3c
a0tBzUMaVTMxdrY1Em7jAy1H4zv952Ql1LHwdNcoi/7cQ/0I59q8fxo+UHnGABOaIxru1xOXl4e7
jrh5m5q1jTrwfaL6AXTuQdAwchHA1A6BJK2sVRS7U5EKFybBhVqc2zRvFapvWT8T51jBV4Mg1XoI
jgsJePkPq3SgtAIIZXSc/9WjQYyI8TbFAJrBDJiaP4lpUfgbjZylpQyigqffkEpi2+WDKZPeXqr2
Tw3nHEbARdvZi3XXXbI6UP09M14lv+mWFmdkmlEIn00a3SZaPis8KwbNHXNLGkGsIL+MG9xFh5FF
l3+GLmf0iss7PSAR+CDb5F3c7BR1IanjnRNFRDewHA6A/50nuM5X1OQhdMoa7f10GWaIWeBweom9
CUFbEnhopTzdFIxzPOwzGe6sBociGhDE3a7tTvxj3o/0QdmlBpemJyTI/xclq4bAHr0d6j3N9DLl
/nHT5RAkaFkSUt+ntdJPpQxpPPZWQ/CJnoo+zXybXkGu9XsG67QOWNIvpRfdL7p5WxAyVQhJKi/d
N8BWEXVEry4B6US2E3YXE2m+eWTCoWYEDgCmCFU3YXIj4Vzk73dDySutOJ1rRBdXzLmZlDhjNAhq
SF0352gcEseUPedxoNyATdqTHOqMr8wI9tS0COKIMjvOusScm4MJpEDaC08r0xSIFHRV7YHM2Gzk
JujZKUeqEnEmac1Tthwp/kkgzOIxkYYkHMCQ41kxr61mcTKEHePU+ajkr1QvsbWX+gsC8LpColPh
iZgLnawF/xEGM2LKVpto5ZyPCVyF1tmooL3yghhTyJ8eta8hp2v1Nu9YaZXesufqt6Js4Zg23YlA
Kx1jKsAKgv3b2Xm63f09Z5n2YA4fg6DDKKfEx8s8C4IOciGiK2wYx5SpdY2Zp86WMRA7RRdoMWpX
muHHDovXE+G9w1ZKWdDFzdTcNfdtdupgi8bTEVCfd4ZbmQkhF/fvsMzfmX0iR7HSz8GfdHq3Sg57
QVpn0Oq2rFy2iJ/L6F8euZT68cRGaNBvcFcezi5Z5D3wV1j6Q9yhYyM18fuJ5qhR7mk0eFjPk6Z/
y0PZBG1gajzgc+TcH30u/WnZdDG/3YtU/7cGNmVV9d18Z5jQ4z6+btX1I/lwsHby5UT4L9spVqDL
WXuPd+zGpCotqfJgtjR8IVZOZUF/HEgWEGHgzdR9OHXCj/azJV/h7XCqi2HFWxmwREya7IvdXdeD
WnlrW8jcpoFjFgl0SXkhbren+zlorLx3xWRQfSbZCfkC4LkF74gqHdjfqV8SK7Gc7XC7Hs77Zmwz
+zfCFsMZa7A4Zc64q+4EwjZt6qDfWHMUNfe/KaP9Bt8Fd5cn6EpMe2sH2z33mppJ85WCF459Kj0k
HknxuRukqqHQZor1MLI0qsw8pJcXC+11Q2J6soEG1Gxl+FRPxadHlgT1ThEZJynxp8dU+z3Ga6Ip
C2T6QcX/kenV81I2yeMKiZ1hrGM0/3e46eyCOhHEcUkHLN776zzxrGMd/vFPFxJmwY8aaZnVn2Xo
CCcAJDriM6ftKBUyDgfzBVbe9PS/2AC2ZG3918VHtXAoupFXzLXUMEnUwcD4KEZoH9oh5V3XfqJR
VKjsX8z8p3qEgwFoLMfrJdFv/5yLSWCi3nmCAsC1CrbnN6Gwg01tGbXZwuqWO9kJLNvKrj6QbuVw
UkDmFRSaSCw0ACApIErhhl7kCk32us6M+8W0b4lGGOAh7LigvuzSSemBvOuGY6twi/0+Ccqw83NY
OCgGx3Cj9jdgXMttkMw3kzGCoc1LjeLC7rtr2WwAO89w4hBQ6DmoAHxExhY38Un7GlrrXENVEGoV
CL3uhVQvJPrLhMhE3Tk0OVFQk57u1NKr7yN4JfpJ7IgD5+Z691J7nPJOvFtNbRpqk3QY9mJBt98e
eI05+CwICP4P9yLvjPg4rIooV0s/9mZWp4TAw2bvScxLXh1G+/M1LqbMKsUi/f57+odssObbJZua
rqhlb3DTW/dXmJ6xcYPkrxkw+0OcO9rHUmiPctlPis+VpJ4Plai/4od3GHXhwzilXoXDmj3AmWde
1xI2zsRRPwxp+bjUwMABjhEH2hWQ3KHNov2MXFD6MMOlwnWm22NZhzwCCyYinjtxjtzAbCteRpWm
Ojercm22BeMiilV3GHKJF/MAcVmjSc5G0MCHXEfmp99nmMOQ6aYViQt5Ql2XxQ5bLvIvt8qgrlML
/RSj8CZ2f/5UWObyTt0U0fJ1Af4sUnVlPET+SqHTwpV+RXGwghadDow6tNZGrkSFhPji+NbzOnm+
N6myo2++3Bj2zt309mScMrEz4vWI9Dq164Q10HrG2s18oTAgwZRu/tD5Rxjd/2nQtYrnjcjfT/fm
qx5odSS5+atHrBF7O874Wh9+6O/crxw1FmsxIvFWdhY1wvPl3MWZHlQk+/z07GikeDO12yZQnrFG
/a0TwNJ6tJaKYQXuD4qsFi8AvXMAV+eZaC4lmbNtj1rh269YITDtSPl4msC1eRd7SnO5t56KxRjr
TloJeJl171KTTijFFbmglqUPJfMKAewkgNeyiiKY8GRmQtxmAZ6wxHNsAWRjMrUqws+xTKQsTBGi
yJ8yd7NRW8gbgUGyNpCM7b6GLzr0Wyu0IOEUQwfHSGCTE6Wq7hboE0aDVyjNM5eZhBnnAZGp0tgg
RsfFOW2CtU/7JHdWpy69ji2k5v7PQcM4QYowG8zMfHNMBDHSlPAONzTvqWrOV8aIr11d38Ucq3Zs
1Am5DW4Ek+QEHTs7/X3g+iA5jeRmhxHXaWloDgXa9gcSiqN+sGPu5hHy0uNJXeooKfHUcMXKfyDS
VJp2A6DA2twsk6OMk62g2W6i1HBli3eUdlOwhQcGn3XtmKQLLkB5zYU5rRnBwSIgoB/0XIFgvrkx
J7nWyPjIh+fD6u3PaJpxMhp0WeuP3TxORT5WIO+xcctrgjF7uteIvNGURSpLsb0/EYMSBGApcXa1
ev+iH8cSmb0V1qwTu9Rq02TnJZt2xsV1Wy6DIhfz2JvD/DMf2/vhvbjQrKJlH4jSVdPNr3+HGrJE
KZT+b1iMIhvg+SFDmZa9AmxiVBM/QQOlovEHReBTS/cV1RMUaMlowh4jXJv3psXMYsbgcvBtUDss
NnEe6DaJ5NAhr1cnOsiD1up/nHA9tZAVE2PONvRxQB45z7cuamTwG48iMrxEDhXcNv9DMlKH4ILU
e9wAK5IBuozxdFr2fWRFctFHIr1Yj8Zs2hXsFL8X3LkUGX5u4mch2zNED3rO306dbzFSZRzBQdk+
cyWYQnzj94TBnm9sks/RUqSjYfGJQyh+F1p2Y/LaqVz/SdKyS7Xp22FrWc0c0+0OIPk8P8NYAAGG
+2S8ixBzqMvDzZCFzlO7aek6AUXBiulXv3fLhy7NajFbSnKefukB66tlejjVSyROmkdz8x+m1z/d
e8HzsKRGZ80UD1uuzvC6y56hl6rPxwYQWUNKcliu6Wi9FlL5OATUt1M060kPLMv7Ct9x5uxmkaAZ
JwKeDty5+fZBGF/4iYxTWWqUPsN+rdvIMG9xF6597mvGIAKNudtpD292+AYSwD6oADZ+gmXs77xX
C6keeUcU6movrQsBe0ele2aNfKJChze4w6uzJRoDueSdbOfLFsZJdAF0oWOKgCt0UkJ5QIV5kk36
s5KUuL1DVCVg0za4R5H7ZhjfdIHkxaLiYVBJ4a+NURUpsgKCCve52UVSgoYUWseAvm0c1t5O0qon
6HEzMpToEX7QvQ1R3qxQEwWaFohY88naI/3XgSXeY+L71W6F9CFzHEKPiovzJeYIjUKhVBuUSpMO
Qg6ajtoHXUmep+E0wKGZxpPrXpG34Qxa5PBOQ2tHn4htpuQG7N8rhPVCNdcDYq9mrzSrVZ0AxXGu
QEdnfOvhnl79PTBf+6YUa4zdk1m9oqK1ZMuaV1pxTvzImKmrIG4vF9Ag5qBJH9rjSzaJmTRvU2yv
AeLY2T6u/QvS4nd2ihLpsIJ4dkeUYRtuKPP59rrwopUbK2vFglW1yHDfSDod4BBiMMZQ/9n9MeHv
DSGxkXUDFse2/OiVypMb/LXYppv6aOh+ZVjwEUbU9E7MqVZi5MAYciymgTn8Uq5FQDPZd3sNRI76
kCm04CYGy8MXqrSWUFEisUbl46rynl9YQl9gqVyBTCpkGF2tooOqUsROb5hVuxJZWPoCE2ouhiwY
/nirZ6LZUJTErH4ONpTf+r0knY4Y88Vr6SrAtyPHZfsAonLbvFsGlo1RHWKY5fXEunuRYbOZ1m3f
BWPSOfMjNRS4Z3+gpZDWt+BKpaanfEEZnFmc31EWd+TcgPFAbl9JsRBdIyvuWAp7AjPFpixMvOBY
wXu4iy+WCZgmBvClL/sopBTiWXn27u9Jw9HMzG79i582uHgN9orfZvfbqeEtKXKRQZJALQnaRH9k
gtvOopU0n/RwKrIlYg7/2OhgGfll8HRucU/KKbh59A5DwUYPczDcjl4mDrPeTYGJWe1Nvm/MOq7P
bxINe7pXQPKWlUA+VA07IgieQqV/aQJTVvk8wZXxNpwW/PGts6tVb4vww+j05TGK0fv0BFyncM4O
sUIu7cmaSjcwdUoKu1Mv5lfapFLlmL3yGc6zZYD8dT6vhv9DSgvtEBWpTkUjYXCNgg35bbrY1Hts
jKusWQVuzEQDZ6JgyvEqIKd1t7iGS8AIKC8FK0/24UbMmnPd6UHl5fc7m4ta77j/U1I6mc9hVydZ
XLp563W5cNPRa4bCazL8liIswpF6afg4gLoRnhCXAOy9eNypA9k14hq84AX7N3/UJwSz40LdgDSA
rH63Ob4sKoVWRgMJHRdONEDpxHxARE4eTQvraQJlq5Hpr//NdJ+Hxd99+0swB2q26/hGXgio7eSO
F+LKf3lmfgC43nScm3gzCw22sT8Ymk3pfVJuPj37jnHaibbyD47l29D2YdZ1qYaBPQpsrpZ9HsgJ
6/7JJ4fMIckaHTCzBBS22qhDkZEFJW6505KqwNSPdwjWxzwyVqXFOnZHEz5x9xjOK6dIPs5OR4s+
BlkOloeuwpn3l0dvtxIZmMX30PuoSBm6T9Bq2L2LzBULR8L1Wh7+sRc6ZNDY1PDHwXyuuM6ToSDS
/UQKnKD54MVxxTXBCOsDB3IW9pHGBM3zZ3CKSe2jR/QZoAueiScHn1BZez5yQLDHNGs9hKstAnW4
n7yLeojT0kegnVjX8ZX2lRO+VArO4n6BAby1gkVQlRTDGpMc6yWEr9LpyGVuYfHMrVA/kgd6W2WQ
+CB1axPoR/AqpMtHJC04Dp7fMzv8z3rhcwl1ED983TvX0f3uBx+Mx7E1M+944t136h515FXPlh8M
RcEOyFGvvyxPmbjlOuug1VXqiHPR1KsS378rZtHUNVxwmK+S5kKJqpRfDVP4kJCbplbd0dKpFZ+N
KkBDeMmOv56umC02BZFQHa05wLa58sPDfk6Au+LwpcJivVCqgUzaP9VzV9wAVwKxBFhEvNgwBolV
I0lQpSr5TyBTKLLIIhiHlHR6F40G+5I7CpXXIp++KX9nZ+CJY/9h3Cf2wcvnMbGxNOu3B9r+KwUV
3o6+sonARqsrCayQpBSznDuJRiemrv7kD56lysgliUOz2ubUN/JhmghjKDj42X8vtg5zqDUjwnMe
l8nxq9bNSbSExIgmdAsFgpb7qxvXTduUfSLoorGMEU9/v0Tnsei6XaVkWsCO+W8+Kq5DvA9c2XLT
P3Rbrx0H4zYzxBLy+WbI1SpukQTASTWgl3ub2iV5bQLlOWmUTxWRcvCgRSqR3ewKvVpWVsO7/kjo
r0qRDmavKxtv4lBtLgxEJ9zV4namF3SW5lUspJMeZ/WRxc1swoGpJcsJGRG7WVPjVQf9Xvj4Y+gG
cS239zbQzqulT5cdZ+benCcJ7NhcHsqGMVlnOY6UX4nGm0D50rK8HXLHu/xaP+sUf8NNxEnElII5
j3G9+Cjl4ASXnETloNRV/DNfQHldo19ze/FC/yWIRin/C31GP12s628qCTgVxKuDADwLTekk8kxu
LMnIXD8MXxYZ2jwmU9ZhwDvr0hHOSzazjdjovaTxQDPVfBrtsJSgQ7hMewGW7jQVFK67IquO2Lsh
uXI1rRMslTgTNLea3e9jX0UiWKV+A6jKjAAbMgGlpjsPKrc6vfIxec84xY/UeSZIDama3q9dqIp2
eu7Qb6nqO3OJce9BOd+EyG+azGPvb4ScyS1sU9YEIkEO+jk7PejKLBHe37FTwCAMm4dHqTDBH5B0
npP5OLQQNbURF5z70X5EsRpMOAbkBrVeYqAgwh7AFKFw8/ZL8q1x/H1ssfTkTNAVZeRQxYpQnJ7H
FKjoDgDDNV9xEoc8SvsZq/8KmlzRhL+/OribBCIyOC2RzEufDKnorDnKa5QwDs8S6SPu3tkKeJTX
CgHOOqlmYLY9cwLz0gQQIlPH/f9Mx+U7KfmtG2w6WP9E+Kbuli3tq5TY3K1uNXHZPQwc5bE/d06V
KbY25k16E8tmku/GJep75x8hQqTQKod8cxbGJly1+FQThjFlO0qeA5V7+0AZE0Xg+28UE3R3rfwK
F0XC+WcvYj0ldxg5lSOQfweeeeai2t5IWjQg8MAL99Bh+eavBc4ok9/DooAdrZ+XPn7Knv2bgjb5
7K3F53p73Wnr1RoTz4r1dVPqPkO+ts6O/lv4SQeR5lGbGpgSQk7aCAdZio/ZlMe9Lw96r9NcebDb
1nLH202BhTfxiF5p8qRINIqY82u40JbnQYTxPC/kM5o3Xl4imgutpieL2uM4g/mk0hZXNz9xWXUx
ONRrw/EDeUgnvHqdUrmDnO23UfJB9HnEP5MMPf+EVUcllP4YkiqSy3ALKTgo6stVv7IR7lNeOBi1
1HGpMviDrk5Hf0quoc/6Vkqfv3QuG1+Sqen/SVBZ9oDkqexURSNweptS1AYbZZvoScxRTqI712H5
At3iXnp7+L95YnRSq2kw3PCUrn63y0WENCSmEveThdoV9SsIT3MBhOdvAmDY9boln8R39ry9U9C5
0uCjffcuv30LNM5S5oiy4TQpzPIu/fyAFZbEKQkNRkQJlmkiTTgCNt0uRPHSiB/NQ96mAQTO9SP2
4TmFgJK2YzQhjJJEcSX2BkLZivRpwjCQKhd9F+hXMo60Zeb1IOdDBE2bSKP13/DGPsWs2VaIrR2U
32cJ+/0wgJvFBV4oXYTD5FWkTcrB3ogocc8IHX6nbvsWB1ui6dmHoYrvWPPcD9O47KYcG9CpmsXp
th57hGudG2kMdIMHl/+HTjVElzuKR2u3lsbD/33hjcieyhejWQne6WUUCthRrrZStCgo9XYZUGcP
bXk/3/zCE+x0clIWYDY3dMauVwLYfaBu90gSPtFcV6ZHhQvGVJeV/+itFDgecJSqy+lUVlVfc+Gm
hjR0og0KX2NACuNwWmr2nUeL/11OH9ebzsPPEYx4+OQGC40BzlFCXwuOYQSzQcYknL4txsHCoh2f
vBTA0Vama+E7kPw2BfTR41zLqMxbyrXWki2weTy4tFIerePmUiwnX2OELfDkGHR+7R/DjYlZ/Igo
MhJqdGvIMWo8rN5uESaI5YXXQdVLocwm1rWijZnXGk8Si1+f43ktutSqa0sQb9nzzBlAWnw3o+E2
ZBanIAIEYFcdg2TbvBHxMhi+6xxXn8cxkyhfzZtnXrxi0a0B5j4QTNWndWA7bkJlMTR/N13zT8wO
rLyvp/dTZJf9pH6vEV/si7NsuPZPvJdX3WWQnq/SYIUfap4c9zvHXl6vWyErowq2kQCq33lv3kmj
HRRy6lo9+ivmV5GySh2jLOUsFRmeFkwDFDQJC8WEbpcgd+Ewlu86yag91mgDpAmUsPBCVifwCLni
8qqVV7THHW8xuLnjLHh9j6679QcA0A2+Qh0erBkpTpznt0v9fJGZpXZt2DORr84ipiTUipeXWXBv
akekxj8EoiXGHK6DHlIMyItS0QP/Cct/68qyxgmBih0l3tJzNHEqrUh1XHvbFzjKxfO6sZxZXJQ9
5NE3bfSWlGs9YEmCImL8EyfKfzSkYa5xL2pzg8tJX7Njsq1VGsgNkjK9hbINTU9eBBVE7ZeOcR++
NTg+TG3UmE6HPT4kZ+Bb8uOHoSZE/t+utF13YXI8VWOaqa9Wh8Nl/52RW3XYPQC26quGSWTb2Psi
H7LCQioODIYqkhCB2RxrUnqCISLc4d87Ib3MO7oud+nTvLu3EVOaJDPHgVjQXhj8YrE9uJ/PDhGr
tnkUjaIyUaPzCXbZqWF9sFxlBBmR8AnE7xwjWt0YrBTjbc9keMjOPsrdzoe5lGMgu5PN+IVpbg7W
mUOUZTIqkBJPmON6wqIiZk9EEn8YcwCiCpE1fVLIQ1H+iio6IKwPfXp8SS9rdK4B31+N/Ij9HBiT
jq4xtD0AVwtSkUHU9FUlCkicOvHKKZ0lf+asbow2cF2GcEcQF/3/wuoLotqjvd7jMMHHxPZE1jXv
t6FKHo0odhNIG5VlA6UZ3WhRpMXKhJtk5ZhsakKjEaNzd/WUWWyA/Y2okTe8EitnleKIK4M4nMCS
oXFk7Eu43WGaH9WqOFJCL2rY99AT60sCp07kfFSE8VGdHyTSA2fFnIxiOyul5KVDTeeEFzSsipOe
8Fx+uZXgSZMimi5rUgxVEX6nep66pnuwKxVpnJ2fUXOElzc5qo+j3Pn85sxiFVwiOTq84mboFnF5
BPuKyUj5GWkRBClOSRASmrx7dE+vv7TVkw26gvqbGN4XNt/kHeOKtbvBSDyrLnhwgdzn6Z9emvnM
9h7Xe22RlBvOpsKGiEk841JeipqUwYsVaMDnuZRiN92O2ILA0pHx2agPERD1rD/18ACZNrLtriwi
7Sp7Z6iblVH36hUcLmHmvW7+sSkH7TtEgjk/+FtqW9duRTptKJu+JyyuDQacs9xXPUp386lvEPI6
Wy1wpP/ernhud1cwfEnngKrs1b2D7h6FsHBRcplpPnjZ9YIvalie+1GFVTz4AV/7FcmL0EgQQ9Po
31Ry0Uly3+dKuKclEPTivelc6mYJ4yygYHm9esd94AGlrhoWZbORiH/z2f2A+nqYTGsxfvtgozma
nb1l5RqFTTVlvy/SvJ8Sat/UjbA0jrxcmYPk+nrgzTjt1v54Fxqp8r8UsJGbkzm7gqNSUo5MDvFv
gk9xvHCc138Av2zBgpq2lYPbTR5PyLINDAqKzdE9HerkUn1tmO9YrFCX/ebmZG0OGVw5OUng1Dz9
ivQZoEkq9wvnnOrh34X34D+4Xz94p+sFLIked8NEOeZTHsU1fqEw+qOGb2LH9VamhPuvDQE9AGqH
IFUGzBLCApBAWAhaVKBCyG6zp/3IFWa1yCYzFU0U/QMtR5Mi5xa1H2SnmECkCJ8/8ZRn5PWTttGn
kOnj+fL6iAOCy5K+f29MYexS5PXWAoHU6LkkhaeNnINnagEWikAtuGW1Vo7UQQG7APmo75wYa8OZ
EdGncKf8ZXg8Nf6Rml7OslKFiqpmW8n5yjHKb9iD0f2+I5R/tpdwwZ93DTTfktUPmijbLvi6PFcv
cwxh9Q0FQI/LSfGANJoGy+nIKie/rhvCJy6/WtlA1Miz0JLH+iU1K2FCGGgQqUmW5hl7U0Gk2rNi
LrrOqb2VSjai/6noAUHiJ+9ucmmhoJeJpA6MV1ZZ8nFCNjwZw2RmiVt50lfskIpRofzD80jMwyHJ
nUl3RSP5wiczwbRZ794k4Y5hOTyeiUfhmt6HlQGhyMz/1nxPd0dHyzhSepR+tQ9MY9aJenYUAif+
EMwXqWzmyTibtS+4w1KXxHhugmV4nrfSfctdF1ihYLH9K11RWGhEgpMepCxDsKUW2jkqPTsrRQ/O
VnLCbPnq92eqh03FUqStqbV0I3EYTynxLkUanstXJ6tLCe6X8LiYYu9RW7MpE4MtauZSfvCYxoaZ
S8NShtfc+UPDjG+oqR9JtxqMSa6QUBR9yqb4iFRZplb4NH+eoC9KW1XgZGQb2wcrZA1pJ8qyr1E+
1uVPEVghWamvRRY0/1Ifia7xIPEWd68p7a706j8GWhwuX4ORrCjktmjV+bc9hhivYFxPCOq5WA/P
HWsi9lsGonBU4UrXoszt+c72E5nXsVBsyEvcYgvfvkJXA7aIXmkqzOL3wOGnrLO6rYWPV2RqBS2j
hz/rGTPBIQvKrHuwBHq5nQ0M/nN7LJnYX0+pzClRbKYeAYbwT0UaTmyPEMVjErH3zHcz8UXT4MZX
yUTlnUdzU0i9hydoxajIc+NX5bRs2l9iAGwnEO3kyBcwbICufHbYPbNZI6Wx9lirJOYA03d+8ROb
SEvwvcsKFQvoxBWARSwHx8zQP0XP08OcoxNKIVNCRII3KQZ1xYuebHBOKcRpXFQAWD713G6fkNo2
zGJVAScBoi5auPbcIhIr0LkwEuxbTutkXqslgkHKhynTanjYC1VjQ8s8JRSecpn5DmGc+20+Fqu0
KwJXdxjIFU49kCtFPckoGTxTu+gX0z1hiaUnP4YGQHLI1jT9WWxaUUwSXDlANBBNm4eH3ovtSNVO
O2+o8q2FdrsgxEOMqneiGgfaG4BtWlSD5DiVHnXRtntFziU/Kfcg9+HHL1DNbuISnK2Z/+qP3BzF
whIhqRFhaBSbvqwZSMqJWDGhzrSp9q+2QZjo/UgeoEMRDCOOnuCBvjTrD6RIABqtJhpDgKI37cTL
I9JyMoXWgpxCggxTGFrrrWEOvY3oSl4HXZjUOVb878Pz7+S75/NM/zvARdZbAaY6SI3PQF72pnO2
rpPpyJeSwuhS6LYzMx78n0L3Hj/N8LiLvC2BZsACf8W1bO7/6u+siYYhjQSvagnl+ctakad1uu/z
yETY7bx2nBLO+SGF4zfwNqV2545rXZ2EyuzEPZyw3IKZvv2bEdUCBVMEvJh4telui0S1q4KwJUW0
mt8zI1pPjGm59X9yl5JTtbSTJvh/ymf4jgsPxDVO7ysL0DAny+20dTmlvtS/Lennl+fHkHBDmbsQ
MmcOhQv+Zy1czm4wZhLun0O5k3kzeKr3qc0BSZDMMN2T/ez4t4m5qnAoXjqjJyGqWDUngmswAz32
8HhqeVVLFfS7vZIx0fOBMm1W8u0AcJAVnFsh9QXI+BdWouBwddYvg3hdPaVqS49JfWkBYqdTcYyn
bY6gpOhI9oU+gCwjP8qH4Y8rNnwJY9UqPoixvEF1396a1QoooUs5F5ldnqKLoFkPMA2wFMhWfGcf
ocoW/Y45C9/tptMj9mqBVPNDszlSDPfx2wsVxQzX+0Du5DWXmmiSVOekKioW1LhjIxG3F47EZ0Wi
LhVY9ZKyveulbEs2S8cLQPtCbVrQXYX1pgDjH98bR2IQN/kCZmv8vSg89ORwKpgMChyjYSPMbGBc
s+BpJl9Ssi2TfWg16k2FXVLAfbeaUjOy5v70+TOmGFXhBVDbVSLtyd49AP/te8dbf1bET3JQPc6s
TI4fo6cxNM4Ct/7v2jSHj8NBpxItBeNCcq+X78dE/7SjaNZV+jOQd9FXJo0AmzenB2T9jjxmFrht
cZq5ySYKE9XciJ5Ra/gzc7y98qqzZ1Jw9Fji1DIdcHg7SEFjQnWFof0u29XS2tBqaFWqz8QvazCb
EKd8XS6yo/wE1Dm2oNUj59wrggMEYxl/SZjwXzgb3sqv80xSKlo4xpVF9UvB4wLV2etIwE+GlJw5
ShmS6Eon+Cy2rfPqMro+wwVaWDSlOHccBbHHBRKRGSdAPXdYtMdLTY9qn4lyg8XvTeMl32WeKNH+
kABjb6qjlOaSYlJsGk8qPTLE6EMQSr8CkVII4SdAQDaF6Fwp2IVA33bgPGohoo9dhaCbb9ff9adi
k8vRI0Ni09LgpRV/LWpWfspQq6mVGHq+gD+J+ji9mqTVpgmEUt/Ogft5fywFfeASPhoqxwNggGao
vNfAMgO19N3+BFnGGlh2s/6UpPMsz0FnTy42n/he183kCOsar0HJR/ROeKL1IszQeRrnwQmhgHvs
ney1RdFSLCFDIY73rZYYbb0O9bYAI43Fgy3rxjGMoSGaZIfXwErMlaw0jniiYRH+UwzjfHbUeYsF
ebNiiHculoNDrSEESnpswNK9/I6Q8328PdX/XkLNgPe3MJmV7Puy1oFxVldDUATYeC7HJ/pEZsv/
Q+SSWUEQL/5Xkps6h26S4Get3je9JfHpElcBv39waMCuhfVLwjXhwRBxfppvw8gQP5BzU3rcCCer
22cQwk0kdnMqZsHbpyHG/ZZxvZo50KR6CBBBYGVg8DTLADdZB4SP4io2yHSah+dlz1/qvewL+g46
xCnpaiEC1D+KlzMy4P4rG07/j4si85AxzOhO6zIl1UVTanPubT+2Sp8Y7HjoU69LnH+aJa/coBfc
+SHEenogFaxoCn6rBp4XLseXEn+h5vAlYxOblQAK+hCeGDDS869JZbGRit8SjBXBS41XHgSlhBNg
WQS3Ft3N+Vit0ABfvFMbHMRs9vMKOM6wySEu9rQ9dkOkvlzpML9GrGWC1BhSD5ytI7t6BuNIWe6d
b+P8K8vYcOrcZVQfFpF6PqVB2LG+GkAsyFKu5LJTeROgsCc8YujYCuL9glb+zz4DuBxBDJuT/tG3
U4i/XYlPImXY8T6rFmomd6OQFvN2tLWQjDhTNUHneiHVsia3ZXdEMfwlqpajASwbuj+cXc2Jk43G
wJ1PXXzXllQUXYvv7NsLDBnkndwQhmxAZoFJ9UGQdi645yKJE+8ax04PqGGjeuu6NSoWobmanJpi
QXzFEjpzU/TXj72dC/uJHJ8mXC7EhSbjDWtyIf9kqizL/MIym2/OxqJa25VMuRkhOq2KQ+elbBWT
/1ncZTYjhERRM0dtr/f0uo6ti0Hp01hGAAp6AJgvXjVmQKhIEUSzyUoRGP2gmulsffwEpYeiGiw2
kDKXAtzY2eYfeEmsMZIHsQ3Xc0xmf/FMO+1/cQYkoAvH7b9jZhLf+wDusghyR+lCLdGqNh5He/qT
/1tH6HR3mxI/uvXk0bg1m3MJA0AYOZMyki/VcFzZdvQu+waUpORKncfO0+aQqf8FI3nM5Rbh5iaR
A8UCEvRM8i8KFynYGRDrYWceBU8o/XwLc4aEndPA8RTz5nSY1Uxl8FXhsv0F2wBkVyr9rOTHsgDr
slx48AMEZdgtt9LDA2+vv7ielp3IAULYRU2QcpYesWR0osgXLX8iMOTDQEYbXoAcS7Hb1moOgBgp
qGfeN24YxX/Y/MpnswFaKft66PCS/fD6l06PtgyvWlF6+iEjeRWM9E3HgnCTkrJ/oQAny0zgz3Dn
aWgyVG7TTjdPVkhTYMVLHGPVajb1YaBVPSFHYs/YrB2SwFYxx1UG3xLUh/ziYITiVygLsam33xJw
E/bsmMKVeIbmT+brGyEAh9Sn0JntMjzP+f9D6+Whvxa0BMjspcTx8XCIow1nUZNWY/KjEQQOMZ9X
abWm8ay9tBN9O6b3XepkgNnheRMU/n2wHS/NHMF6iCqixJjVqCv0xe+Z8yQbZZBpcTD5C9I5/uTf
Wp8Ir5/gnQqbfXo3myNSMIn4Oy+0gPU865bzxmGZR3iW9l6WeBlKUAEm4c7PmcEltlk2Yj5c6XZK
ac0i+RdFzFI8DRJhlFTa+Rubhk8SxUUWYIVbTuPMrxz/BhSwhF/k98XtbDjRdlJ3Ckh9/2SZ/Lhw
vmVP5U6d0ZJf7W8HPTtL2OfOCe/MIKPohREVY19YdLaTEJ4XZ/flQnQT+e47QRdPS0Cqxp6AtKUO
QDfUgTnoZAQ1IHiLO4U20sE8CN7hNQFOnLML6slftpWxTJIuEPWoP6VOfBWNJ297MC9KAgtjMMAl
kNNJI+m7IN0bpOCjhBdknNDo9XJCHRcS5ZatipojjiFcHVQn7YDCwx5Do2XysL8c1soZWxZQAzQp
RWUNZoJ2Q6Po4ZzvsK9rcxm0eIw0gfm11mN8NFOLTIXLJW22ouAFsQIo07DVGpGbkzY2RDyv5eY2
DwrdLsbZOpSO4/dUrW9y4ghCLy2G8RPskVGiDQjJQKjWNl7bDS2PpzywwEfzDAv7RtWM1t97Rbf+
WlJu932fOtR1aio8it+CotwWMbJUu9zR9F2QGd+YjQKZny8FwJQc8z9Y8gGs7nRKtVvNcdQrJM5m
MEtWU5Gxn5y5d1yA0p+uBsVEV/Wi5W1n9juKDulhxCdKiDoNdTrk5ogj++iyV5zpi5fmoc01rLPs
nIpQBMWzEw6OymO+AUgJKnkyFSXXuX8e2/fDcQ07ldUlZhLTv+6IMehlQvfXTArlnz0wpVVFqefP
3+04lfwBLOBG+byT01gpzkfo9R5LG8eqlvgemcE3phJP5kkluEIp6SlVmUGqfJjnwlq+h3+KML5Q
m6Exqx6UDye+R+W2OlfOjpsVY4PzZXbH5NSGvHBqOv2/NRrbYbkQvPd2wH1MVLc4nknkR367GmFG
FN+Q83zX1NXlFA97mAsxxNGQVxHMFKvUwgkGVoPQpigXWjf5d110nIcuZcXthrZhAZXtUrJrIJjH
ZDIPKz6IWMnLHNfRiqUNF+Kp6id5wlCBzukrN+s5OaPc2NbxgSRLOzMFpwa+AMZxbC53BgZ71p++
0o0YJ5FYftPf9/iaeNLkBQzTh+n0aPUB6+KI55MDvOf3WRLBJcEXp8AdVawUt25v56eBlGILj4Qb
hVtyxPnYsBrPMi1/uYoHGwGT2HgR2M3KJLTsFPgHt+9GQDp3gFu9XJU+T/4+AEYiidLXGC1qXp3p
G7WQWFVaj4wJDvcGS1z9UwiuMFxUp1cw//OvikNyEX4ZQ9xbvTKgSEhr7c0dtRD4z36UwM+sK0h+
5PYvxA+ZoIYzT/EaCnLZGBcqI/BvThkPlMT129+DDdDOegTOddHl81sknEY1GH92rd6JMli73djz
wHjzfkEiAg0YffmJjTOfKSwNk0TqOQkwY/eJFhN/uir5eYDaxmvQLL+Mnp6zPxQTl0OqrGrHzuk0
mIXTpTojAyvxUpLErmlFGdSfAQI2RFFQf6WPxoV9F9jMZhdceDnbPulm7i0Ov+OM0T2EnMzuVtli
pbZMMPlhEFPN4hlzaXiC4K4u4DjgK9tl4sygan+5/bgEIeu7pWKkuZvzJ4h+clbvUEsp/mC7i0SJ
mZz8h/HZR4mOQBBqHdNphAf5E4Yll2rWq49u06/uA7cPT6lIA/3pqYEthvSgqDwjgdc1h8qnkuLt
4xrzuzIgeiSpLAgPW3Dx/LBnM7Qy95NrqrsBaUUc4tmFBT4spIpkvtb/+TTXEYcDm3RsmyHw5uxm
ky7Hp4FbcDKCQT5PXhuTbPvkOkCQYVvB1ylGIpN6GiH4/mRJeae8c7QbM/Iq3DUKWxpc//rDm2mh
R7BokTuG6uCk8dIMOAJO8pEAklUzfrIfM1uckr6CY0XWfitCeVF3f3+M1uN6o5ya4zlpWoc4fH1C
BBYizK3nmludH6nxopGYwaR/9inRhKEfIEj9fFZqRpp1Hm3dxlOqtFsiXUzeCQNmVpAiuJ6nAoWd
mVBBVjhhV3fz0513axOzNrQSIQhr+MEPWQkXpYI1cLjLdBkgJaXrUPW/umesYgh9rz44eLon8OVv
hjo6lL77QfwfljJ0tAgXI7vtvN8gkTaJi8tcjWI7RQdKalGPA5pVapudRE0Y9jrHNFXBjtF2pQUo
mPG7uSgnYcXTuw86SrgKJ71uHIxbVMnRojgr7E0X62sn6d5oQ6APXkfkgKtxtBA1wzEYFCgcf37n
gXM6RggXrFM8MuZYDAitvDX0rFWFM97P8JA96NISNNnbk7kq0MFUUJTbKKcGb9cQpAfBEyHR/QcR
Twfu+Z++GI/wYPmeTo/KvQ+v9NK2DEV9X/n+pI/t5eOe/dFovc+b9AZ7cs3FtcqLncPZhjyqnmAK
ARTa5W6XRwV2ejK7aQdU95AqZQOMAA7OOwYSCR19mHH1xsU8PFCmYN78DZVlKX8f91kcWUakfj7p
BjvVJHjAPo7SX3dw58/bEPqzGqPu9kcwdNTHIRkjGuT3ZoHQsMY83SsLJOguPGLjID3CQYNYOB30
E0cB3RxUXDfl3W/Wp717DV2a0Z0j2ngzJu3T9GrWvfkWOHEJ/pLtljfC9QrjxFBqX/zS3T7eJ+n+
iDJRCA154x0gL4Jn87eZL3KacskPOFTAdJAUBPK8U42K5kMQ1nxF/PNr7exp45tcopG3703Ab4mZ
bKV1LKi+mlK5kDcqyLBvvXNjuLs3I372/G1K2WHnUCQgFCM05rOR6Cd1EiaZhFjUV+Ue88Pm9mDd
e6vxwxyb/UInNIY57hyYqwFNcy5xUAQNVx3Cf0uN/+4yA4pL4ck7zxPndaYD9MeT6wRmoIFTvMMb
j6SBSLsgehq3YXLunxvKu3IHK31DSIuXthWsc/9tQE/0dZszsd1KD0yQCtCIg6hLia8gDcJsCmw3
8W1Xi8yvjglC5nXvKGx2x+OkYs3m4gvaPRauWXgRknFyCkEXWqXoxI8G0Hq6x64hwbA7D9yXCP/h
vHgR/4zLJ9bp0F1HXHbwNYS1h5rHQJOTjaTTUBytyjVG2+DKt2XTfdROEEDAnjn42/GLCHGYh3Ii
0eQLx8QqZL7vlLNdzIrVoLHu+EIZC1qnrvDLJmQj8JOHqorRLjO8Srok3aoMN7ML+EA256xgZxbd
7lxEMqS6DBUKtvP4iAniGl0CSKubOirxbSOTJZ+HnPHAxb6C42fz/rR0vRPbT00sbLE+YLT+1HKm
75mVatmmPVhrdYXpyISkTYII/Ebxhvo00xBMcIln0G8bwKZaYovxO9JWpT7LW45tIBffvmRdolxo
QiZoFIriZgDjSo+TWqcWNKFTvPCEOO6jXKot5mDcLUet8oFTyhBh4ujkq8IUCNhbZNKO+vfgpnSj
Q1Y2GwD/1RIsBLphDguTDWcnPTs0X/b6IFzxEQVaQg/Ke7eInD0r5NJpHlR+27ZLhGQsrAH+G+YT
2SUl0HFSFjmsu3chXHPOv1o2gU+1iTa2kT+hqParLBG1/B2EwIUT4Hs8VTSLiw6UDOVdgaS7bVwp
SL7/2+lpeHVjDQsFUXz7HJbSwyu9cvm+DsXNK2ysQUW1rhKov4iCcgRTjP6JY+05ptFF3Ubn1u2g
1mDvc24urAxDUmiPgeSbjzPuNe48CTDL0HeSj8Uljby4ys35lfpZlzlP2YZGQgI1eEr6bZLdo6B4
A5cZnro0x8TgUI3573KYSO+Kca6bvpuL7VHDurbZfWFLoPcUT+0/WESbXL7ZKVNO7IbA6Hf+MUOG
larOang68GACRg+lDzgkJC6xeGM/+05QThzlvc3SrwGgWoR5DmbuLeyDRoivklLHyk3tdXs6CgZY
dSfPpQTM/MK481Fqh43ffCaSr7MKHnqJI3+jIZ0fx/zYOkxEYpKfO1fE46DBtQCEU1S7peALvzkl
CLl2Q5MIs0O6eiPjJS0tsmcst06pTY2TErvZrJTJzynaEqf8DhWus3nm0Rt7ngYdFezXPEoI57uI
s8vdOImy61HOZehti2MBGAtqYWGV6KsZRlGutfnLYfM8OdNqxSEqAiRpeWQWjEsHD6NJ5w5UGKK1
6cFfXAaDrUhrKzol/mj4+tN9aYGEfW3AUzMYcUwIiomRWEzDbC4NfyKPWOYilvUv8PVdVLmBqYqV
C+AHK5BB2Xuu2j0rKkh3CF6A+bG0NBxbe8hdSwU+Evyh3gSqNocbV7TDpSRLvNxw+RDgKkh8x8MG
H1+w0H1nG08w62cz1YpSr+y5TlfOr/+akvF/+M8MaVdUZUs499oomEUqfdknmIvpSMq6Q3ocE7mc
w685AlXg5ACkrQnC8OdKbxHoMYwcXslzsLRrkpXk7Ezn8B1SKvxV/dGi06qE+M17uxR7IYwhxb/8
fZD+BmcE4P1rpfi9fuPeaBhWopBY6ZKXtwUmGOiFf5AfAMQ95dhXnqYrZRlLVW6fvRCvFQGwrKNY
f5qN8qmRdMFZ8FBv1BFsDL2y5cDPN4FL4mxgp6VqqmQMNrDhxB7Rn9CjZra3/4cNTTl8prMFraPj
5Ug+Jr7WiPdNa62EM3r4ycFT+Ts4Fbj5ShWN+2giF+3ny7ns77+QHSiJhgFWn+kfm4+l1KdPdBNG
fyA2+1E/NFASRZKKFNWdzrseCmES7J0hS8u7U8w4TWEuqb62IlajWu4KcV1umSLs+6l5XAzZ0b3H
k/MQ8LlxvSLlRHEQUDcI5o8pNRbFbk4KsVtaBtaK6vS2NpgnDn1juBx3rS8coO8usMEOukYDC7YL
tnEQEwHvjR4teu4OTfUXEXbNptXXgL6iiuCLgL/YCJkZf04G/gj0Fkv4Y+l9j6BWKG/Xt1U9h57Z
gons4YSvJLxV7UqlBpzAEfRebcFh9E8jFDUxwc2hZumCTnBHzvTgpZMTBEdm8Wo/G76dw8rMIVQ4
W8Y2872PJj8XqdaBHTFJuiXTeAIB0ItulWn1HDcWt08ysyFm68cHYm0K+mWrsZxVQUXAKwUycqQB
ApMkOXXWnvSUwONIv+ZNDpjb3Y1kLcTaL6hMnUUE1lwACeXfm5TSGrr4MNCpUFwsL7tFWMmaUwhY
pA1Xj17QqKnx5LMK1kWJGOhIfLORdieL/qoQl1QdPW6l6xG2tUjMkMuYflq1QR2o0DXyA35deVaa
IzvjUQQTzwjrDIy48OCGkaw6+AsIQhjvpMOscwe4cNre4b7qXTjcU7tVl3glQFHPAgjgXmEuZAUo
JxhLbhyOT/fIulHGdjn3CDcfncSErMxgdhT4DXgDLz1PCn8sadyIijFyv0oX99Yl13NbuTecMbgo
TeapJB5EemmjmJM/Yzx1JHXHjClj/0v9vRgvY/p0r4WJNUkIgNKfNXhTVAmPag3Ncr+UoyCAI20U
vi8YqR06PgxrG5FQ6ZpOi03wSe8eSS1oGSlGNwtIgqwXyITjnCDh8iXDVZRF6bQvJ3pKUe2pCq2x
8kgo4MV6iy0XhGDkG+ywn5+l0+wXEX0Ud8dUiH3NPf/3B60OeLzqf2ygTQKvze+PpzclWMl0VO8B
A3WQ2GRLACIlNVawEoRP5YhiCRXD00AMEU48l8C3d991Cc6u+OR0KyEnu/BlabnEKyKn4AyrRkUA
uGm6HKwUD1Qg2ahVpgZso4UzSLkDnB0VPbYsF6WaijCZFMeiUO3KK7gmCDYmh0e11cf15SsCUiN6
52pC+j9eqTlvMQE74tD1EqBGQX1ZJIiMOHPmDElWx+sOY5DapDi5vkt/G0vAgQS/Zi+Ku8Oie7x5
MDWhKyFrDrdlsrqdsxqCQrB2Fb15CXYpsxZ/vmelWUzJikyXZIpnUx29+wmbcRZ5U7y5eApRh55d
JQaiDU0y90efWo3wbXBZ+TwMucPge81ZE7fpZricPuKAOlvDJjdcuImbLVWxTAJSu5rTozp9PgNe
qSYlRPUrqHLhr8eurKzoOjctr1uPgRhwIHf+HXFsd+t/nh/lBLCYK9oDst+pnCB6k6eWrD+Q6jc8
Fwxi9YkxdP98MxKQfXolm9yuzKbMihAPwFQ1IXDxSUhzYC30ZO+MQEIrLfn1YrNpzpxSxYCe9p8l
dSq0eQZOgSBuxBBqfF18S/LyVQUckpM/1hlckxEcABk3GIH6hD3OmJBz/F7xc+Xj9G4GBrVlyDav
2srRMPYCA8t2Tf3Bzd3nPc4tkv038czyxsq3lsvRY5Sf1DZa8UbCTl0VB3lOI3QMcwnuQSuqJXk9
3C+hOpA54HpeyxGy6p5BUATOk6PqyTbpHsx65Sj2CqkiTAvajZHRX3Sm8ZWb1UXpryGQH+y9Q3fH
LSZ4zlxf8dhkAVBhdCJJA0C4E4kHIEEtLFQcTO1Zvl9QP/ywLpnYbKeOdunNlPx/GzPza/7aImNb
hzDW9Bm92upsffWQfapW5709xWejGKJWgEeYq47dlnK48J/k66kxhuJZSgaumP0oe+28KBebh4ge
WerBd6sldJ6i+CVhBb6psjIOVbtit74uB49LnqAbY4ATOL+Af2Pt/VxnamyZ3mGSqeeRfpzPKUcM
ABzsuyg5TbHUiuI5iVQKiHixBMaGxGcK8UfgyFuNvMuGRSHnHECDqnWq+eAVwBDM1qB8qmeDuu04
PKzfKEXcp+T7nHVEWa1zcH2aWm9XkIzNx2PCkwDJ2GvSSgFsGVQNgaKKVbCnXkSpOTEVRIWwSJ05
1TIpEHbRH/Q8joIqt9s693YvRrqv13upOyuMMxq0a0NFvifJLXEAIkE3GNrcaFgZOhbHwHKyLNOD
qi9h0gv8RDkpXXcfq8maWpA9KvRJW6E+IQNOEf5vUtaXxz+boGjp1rartWIWxoboJXeGEs1vzwhM
Vkcvdfu7ZkeE97zz0QSI2V4rL4mQeMXbF+NACPX/i3RDd3yZxGnGaTTp8sPF+h+7O6AAK/hm0LhN
lhVIQEH8UVIvjdNKlDs6W/juHVjG9P5v9DfpKX/lWUg7B7BBsp/0/wlCYCMvujWY8lrWvZ+herxq
FLBENnAvKnRHOhXawVk8X2LLOPEOH7L6NKJzdhPJ+rgvfkoRN+7bY7OVhXVTChJ22nAXkyw9NYQE
MT923Ian4WMgeYpn8KyRf1qAWLAgFtTbxsymTFWz0akcH7lhacRN+ZLuW2DkvA84t03/9jo7R4Wd
BuC29SeMlFvpOWVZC3DhNPo1e7qv65TXQxKDeWzjq72zLZz5+iqg4Dqq+lgyX9SkrhC7sZnrVJzh
BF1aWZlzd20eOgSMSOH1E+Lob1n88iMFtt3nq43fKxIZVeZGgl6URT1LSkGLfr5aA5Q5cjG+73jV
mGEPlWxvfIrxcOnWp4ovYcUsn6lUG6RwEwYOkWH8fx4F/15Z65//qW2BEWuJetCWMW/EF1dz2S8e
Ru29vIf7YgyJWeDJUTD2jDi6kjriD+2h/NkSEvr6iKaYlRi7ESouGtX2xSyDf5b25qyUr/D1VF67
zVLx5gWaqsiOHRejNDlqDQ5CW+7ogEJ72kdxGb1m2xnd6Lj2A8v0GV3o7nCUVkldNOqvUSPV9c85
OLBburEBdi+acbhs8ifQG/BKVI0/CZmxV2FN8ka2TzQmqef700uOpgDSKBVAc3GUeX3IApiT1Mi2
6LIbgcExj73xPetvNL0JJX8YBrt5tWRaxDRrpLHaqqMHV/5kRORL2vQdUUWaBYvnhUOPZEPl6xKt
LoUX8OKkQLQC1IU7Aub/89PCec0IrV4cEAgyqQd7GToGR0fC2+MsPPyjA0SAlvjPgdrK9qqyAFiT
OtWVblQrBHVEyE8PdbxCjrScs7t7rXcvCzIlskd7sIq939k58mJi/sIBMohh76Oy4RjSWDoXawGX
TnUQaR9CJ3wht5bDOoy3w1EHnoR14Si5cAZIUBWT4ThHbqbHI+QogOO7mrWe4Ac+VyBRhFkcbaxc
YPJ8m4s79mul/bI22is0v7DZWiV3x0hqu8ETJUT886x46a2lrFt5Icr6larwKGcX2OHB0vta02BB
LPQT7A18mjDQt48aTVm0CyoeeyqYtYn1G3SdJy3HjfjxgZqQDdBC9zo9x7qH0rnPWXUZA3eBSZBX
gx2WA+9/GCJaq94DceiIxzQn+M+n5R2aLNGyLJaRVa0RsTfirtpmfLY5Rkpro2c+VTl9F9ZKLp+p
PmLYHzt5c5hmkEUwAtWWoZWxS7BkIetsoFVro+E8rWPC/and21ylZk0o8IVQg850K7eNqzxF8VOu
vciJfOmKIb1b/0xxRC1/bFB8IffzTbsoTTisTYjtOhxITQIGPXdArAkI6TDVhfdlfY8AhgO7Hf+S
u3KdG9XChHH0Zc+Vi0Sztpqk9aT38DxpuSVEcwvI4RmSNbvfx7CBxRl2nxzXPN9GAyg4eQ1OIPR3
9arDpXdsgIVKLdTgDo4U9chKJd5OdMBgQ20y0bbsa2hbbdguRjwiQNa6qx09mwe56Y5a15lshr9S
oJe7vLnTgb1M/xDTx/fBywDjbdiVN+jJ6DwiMjWqak644Whdf9b0xcwSaEJjpKdtodo2EP8UzTSF
kqVCg22Q53EHwsEyr8ZpK9aiiYuKtdhZlnrpzi/kPqA8HD0Maos8lpypDyTQPqJ0Nv9DtTjyiiWp
EudODk8Dk0xAu43dcF1vfeO71LUgxNEsUcng4eO3SCAnt1ZY2JxyXNI6DaU3TD0z+VmFOmmet90E
uD53MKSD4NXfGMb1XwrMqDGIGcmYpAgu9Pqr0BLiTFqC3nQI7mXGIQ7S6ZhnfgeGfIb8aOF9EtCR
BhLMsXQLOYxGr6NjzQtGRF25yVDy4fGm6DiNitaEs+b2GZPfFax8C1CdLCgRT4qq20nPebk5uL3h
VtPzZnzhnZECGrVriszx3hPG2UmZOlyr8kqsU+Qwf2T20VpT2N3tlpWP6c/UA/2THWDRhXuFcjaA
fuO+Tcw6TPXssm8hsCe2lR10CuKitQIJLWTiEqYRrpK3yv/9LMff7E4rc4JNjQCBpda61e39Cfx2
nlyHYqYT+xms8reQg6n+idYOFCJYb6eEU6PYpjG9AL5YVphcJWD53nLKQtosiF1FI8Fc+VYbRqoJ
EiB8gvtp4LMHPWW6sR9VSGIxv4h1ui8N2TRdK7yEOYo+WM9lGHn1txV2TtX7Boh0uVs4YSBNeHtY
uZR93rosC7RehO8oYyOqZTuJFPYSX38JyY96tKbfUo6yd/63pbWT2uxIbDpa+QQdX4CE1QvWczPj
s7s7dLeBDmU0ihtYbpr8pFMvTz4NAy2A7+tZq/SOB+yXwPVkSql+cceQxdnco84LoNzoLnoAQ4AM
8aqvMD0IQrTU3KGmqTvxJRqX8QEGQO1PXwELHHYLlWz7YtiWTC8yiP7IDqK7onORxRYMHIJiaBhy
Gq6SQZ5BybN+RQkOeiQpt7axw/X4RM79eyiEPIWufFzcc4CATNMJ0i/XIiu3ttyq3yy0g/18AEsV
R4hoAMisRqlERpJZaQqahDgqCfoOy2kiU0VJ3YG3nSSnSKTdqhLKbaQyctVnUuhWXDn2MNvZyOne
Xl05VeqZ4JvzFeNNY6i3OzVxisbYT0nOSqlLAug05aP2y02/Wc9qMoKKKtbWz5Cx+pMiwYVqTtdn
p3F4uyTGVP+Cegk3uzupSkP4Qxp26qioVR4j4B+gTV4ew048Kmze/arPcxE0X2XB9GNeeFL79Ak5
F+kRWOt57JkXSEwqwc6NLX+3/mrPUOAd2o+EJB8DznZ+G/upgd+/dUa/lhSlA6R/uw2OURLUQBPH
+DyPAVfulm2+veUOwm/W+lXix450GSVkHOj8zGnMp72q78UUg9LlzH5dO251k//gMhvPAhjCoE8e
/I8NJTEEKlsOr3YJ/7Boi4PvrTPhTCK1a1BtSF3CQ5k2uz3MmTR6J0FHSNHzrFkiEqjkJAyB7z+S
orCgEUlLZ9YYDdQnDzjPcZ0PNKF2re9zlVHvmJ/fu/RitZLof95vGleP0EGpg2clGkrK/ksGTR2N
KMHQP6wNyKLZwZawTmwi4xUFftAiT+SFc6RgZs2G1n8vPFmVmrzWd0pExgXQzxWQwo4UOhdWA4ek
JGGH9f0D/Rph1al2Z0/u33EF6LMokcjp+605LOtaxjV8J+R/AJQ4oJ7p5oDO1F3322PlmTFfnMAd
NyBBL8WhGpfhCOPlUXMszyJwXlhGe2QLHoLEzfGstxY6XrEDKgSdDknj4M8G1988+G3M3RAeszrC
m3S22x9rGu5SQLnRFMaFEwydqAyd3pw+MXECcuQ4wQgtwKBdgjwyEIYz5zE8W8yBdUn22SYb5PC2
QredT7VaQ00kTsDxaFQL9FNG60PDSMnI7hr2zTPsv7U6VN8XlQQOaHNjGmONRKg2qN+IeAYFtVc1
YSoR8V1fYsgqt5ldt18TCyqFEBv951Rx0eqnCZBvxiNyZSZLMqMXxc6IeVd10TmMehN1lrnYvjzY
Rn5KC2t62hVaie+QSQhM/hAY4Iwf4PeUxNTVyoHlWK5EK2ivHzOG61VBhsZLdY3FoWiVsHfvvJmX
MNZ05Mu+fXy/JgkzvkFmIj1HIobfGbYmsqeJj8uKopkFQKkuOl3uJesqw8Mff+Okpw18glMaU8hG
FqtJ3fyHVOZjmtzZwQz6pH+KJX08twosjoPTyvoJ9wW+SiWCP8rfgzp8SIKkJ4R6/52CgDCoTzPV
mxUXM6ougjLhwsK5OyBm5vAUYq9NXHewcDG03LcErGVL0YOk/FyesIZxyxfD1hBacKl0KCB3tcwA
4yGMoN5OIjvzKSsHwpiyHDo4wz7Rd28FfGxHLPl4DmYbO08cGdM3ATbCbxc3wKg4nzJHgyZmHQo/
Z96lNdm+YMakZeFJHauPKOgfIERxJvf2n2AwQtJjNni39YggxFyZQ5fd6s21pV4OVO0OPNrzf7qw
zrVSW6dOBT/l24NRzhTjbpGpHEkn1W6Y5iHEujDpYWosZarTgqTCxz0Tk1/et/yAkWmP0tZ5f/Fn
d+suzkAwF7LPO1V0d5sOrvVYr4mvcJNbJ/2jpUW/uSndmjFVdpWXvKKTRfZY0di7hH6SysixgFOk
SlMWWLbpqU+QNa6biWyLjJ+v7hoH1c/T0G/Z+cNYji2+3xNTO+hmh407PypjdWaYCcnCtgNAaFJx
gOvzFQ8F+zzYH7wjF1oqoOo/l1uAi4gtaKQuUBXNbwMmfRHOxRU7swHev6DhtzFlRNC4B7Sg3z+j
Ffw5C6r21j+eV8OYsnyKxyb+B5CA0LiqM778dlx+FvhGmNm07dD/eE6SRLBvFiHB7PUjkeCOq2k8
ol/12i9KJpKljNcigz2ipfYm5dTsZI8pcYmhLSMKKNs+DGnlHvQLtX8f7vMMhhE8I6UJYMAeox4/
AXcXmMG5y6ceGmMkcaoe6K7rkaMffKEbPhbrjpnlkmtUlXlP2gMncq1MZEY8TJmkPSrw9xauVdAh
1lwmIbzJkaePkaCDDEtAXiNEKnDwLSqx2eYTXnzbvMUT3XhxVu2ekn1XwEipprLcKQmtbQ4bvN0x
hcFISMXdZaZSXoe4qJNUzZ5OqfOBv2qTEHEBXKLGEF212IBloh1XBJ8JLIEn7ceUKIyT5/K3O11i
WeA4n974QYsaFNzNbLYM3Gj+3qVb1I/i2UU2jCehci8xhjJSENuL8HRkEgi0R147j4JaewR4dBQT
2bi1VoeyDxKNA12qv+zPs1EugAiyhxEFqvFv065DoQM4BlrOFr+zV3343tX6c/WPrsihxFlxqMrq
naYEa1mOG1+wiGMQ8bMy5QYaEBkF9qK5KfIztoL3qc7U75VzyHFDcsuJZ9+un87WKcYmPYH0LPtP
JiUdDBG8fM5gOhBI6s3wtRPCfLF/bGnRhoItw995gsWLLG4mbNU6oflKiXNg1WSAQNGVGwFE8OUj
KkhFpawb2AfFczYSJih/aYNZSSl8/1voA9vylp8HZ7NBXbirBiggiamlkoEfLzVCmvt8/1C7qnh9
uJzZFhz6N1nSVTyf3pORqRDTQCdJ5X3viQELtTy1oBsEAZO+OJV/j/DfnL1b9/VVf7ERqttMQ/sK
yYexSrV+iGsN2wZIEhiTJXeArDTaUVnltTCUlqrPMkl2qVpwKWAuf83TDpku+wIgidyyJWHkbmJH
FL5tKYXC9+MZbsw8eBj9IKPMJKXEcCE9TWwiJm75MwB4rjFHZaLsrHrmJLd2sAz4TjGRZAkwcr7I
GZhYvbYsfGcwmWP8U44FS2DfzdUsCj7H+sSZ/wwRGCLeSuChQDZahosDmb09nWhlqveG6QPKX2Sv
eDyYvKBW3ybrt1iZibpGH0FRFWOB4i6TQWPB9a+WLDfBHOx4Zc78Lvc0Zp/zL2T7tecds+fXGp9F
o7Fin2MbqY+fahcrO7oqLP4NhtWSTJ9N0h/fF7AFq4vyjFVPkqdFA/8DWjsq0ou9sZh0Q9IqMrOJ
SDyyiNganzTylqTreIEQGOvE3FIOS+cwlA7NOr03aRfyudj+288BsZfv7QforG7hZ09B7D/Fxbt/
jFaePsmfBv2bBp2gN0ztEmOrCNEnMKG+o7a36pIeqAv6KG4NIFcm9aTpEydBt2mtAeUAGOKF03PH
JJnlFY32hu1THlbgv6ruILFcku191ue8yy02RgmT2bAKpmZ/1KRlZxHzT/rzmiFb0nHSVCSjMvke
sPZE80lFtGd4mGn2NvHZdZD45tWer4g4yAnRqU6AIBJ25C7hA9TUU7MYfOGbI4LgUHlFjFZP15A/
HNyJ2DbBMzJ0MYv3CEg06xnl5aScTaufeGknfyGZyFFTqcb4rz1J2n5XlzZE3Mic1E2RwuwMDFwG
ramQnvfWudXP6pTYQZ95jLLZPmWzZiNYLKeEyfZ3heOZyqBKMOjlSxZUEwHknOXKRd2BUHk8+NOF
1fOqw9+v6ZibChMPGj20rUohvYLozzJ1BfWtbNLyvsTW0UVpqggOEkk9ibufL4nqcnJjU+2nuduy
SJsDh4354uu8alRB0yjLVV9GBGzM5+bHOiElJh5Cudn/R7S8xnjcQviaYDrhDUCt1QJ5oiu5MVeH
M2Tpys92HnbFbv4X9FTQ6rp9MIp5WcLbYbpALRSf2GeNuk3E1h3j2RVr+Xm05qrVI0Hzfk/T5k59
oFWTUdNPslegMX7ZuaVXT4QkP1vnK2mEzCTG/WKUkbzrL6YP1313GVZTa06PslJGZclb+pVC4xLS
HzK4nSRpuiTdoQAXUpQluqi97cp3L7j1KXQo1A5iMAh6a+ZswL521mmsVmHTuV3rYrmVIbHwO4qS
0pwGATzYWL3kz5kJ+0JPURf4lhqfY5yxJGzV8ref3x8VsszabJrJpq5u8ggg2XGADS8lVG+DD1Sb
rDVx9u7chiAvlLygLr38pCesyiCjDreZIOUsiDJbOoVE+4FnnewaDJK/8ZBH+lpFDB5mK3d4mDcl
+RYoIsbgNzx4n+NLZ6kLLPLoMRoOho5dKU3u5r41I16RrxwZbqpzwo+8O5TGAEdbqm1Vbq8cIpOH
T3nyWDcB1NXUlZlu/0iC5p7GzV7jMCxJjvy4/Ui/jZizwlJRbGBHdiOg+QLOfkF/K3TI+cF2S9G2
evoupTTpvLv1+vmsLxIoNuzksq3wpfRcoz6aRf88gjeCLRjutLYpvB32uup1pFwD1654mlFdVxvV
E6XuZRMP5ilZb/qq5uvsOmKgbHZH7CSduMPJQXtPVV0Ine1OdTeB2t5PTjhiAXej2MbEUG7JWapP
suPHSmGLGC8oQFmIVkCeugvhK63DULwvPOnH/9iKqDhpJXbvTy5PeoGPyQPZrAsfpDcePnwzE47L
xHj5lgj9mmTaPbl1w8k6O3Xh6sk2g+f5hHe15v18BcWWFB6HedE+39uQDM2ZeRG7kLBWmB7HVFs+
xG8Ybj/xUS0Zs9oWRby2G1p4gTVThlEj8iIaSyQ8t47d9W+uSx9ZWiLPFkOljnFGIqg934lfODXC
Y40ZJfPP/+NsEtRYfuErunv+vVyyzmH+U4PdqPnLI3SUpyPAfTa1CaCPxbrptOFk0Hl/lL8/kN9h
VBJ/soYszDlbw8TTYyr+io67JE3V4aia6Ql33NNgXjJY6JtKf+sNSSaXZ1hP0IR2sz60iwKp9HDJ
AAyYZVLa76UVkXaVgr8R9VBbXdPP7cUatQV7G/sX5hIlxCBVepeNZ42EL7hh2rEWrQjMGTCQV569
9Qo6z+EJkXVbWPjSHkCSQwVCZemAHJNzLCXmpgTaIldMLOhMyQYi+OblOQ8CwE+XXTBzaEbzyQil
8W+MmL3cOmYeqr5NQKdGVyoRXFwiieRZDZq+bgXAarMcMpVf+wqxLMqFzcA3UyTFTyHbXY38m2Ot
9zpnQ7PuZ9pcJOr61EG/TaE4Pm6MdiIvsN1kQVA8rIrb/bzdIjXKklkvJ6EoroNJ14iqqolMW824
4/nwX5dVfm+wzI9ePczgw8ogt3O+3INU/MDg0bX/Lcm2Y3SuyFjxUQblakjiRJKS67MxBVycUpqU
I3DM4d//EgEz3ClB8y9GIfMM7Na8oasCbHR6CXkpzJ7Yo0Li9FvTboHhU0QvwGDTzWNtBVuGgEsV
ddpnBI5smE+f54GiYOrhHitZh5U5MJoBLWOKTYUOfcDQl8oqar3/GIK4bu9XFGs27Xp/BfF4jsTb
HqtpzwHioTZiSlHW4bmFg5NQpy5OgN16xDoFjT/yiUNP8Sya2okUiDnusWaigDzDthXrlfMgrU+I
xibCcKNyToV7/F4zmy29T0+Lyb6TM5TVJGB0UL3DTsrO7omrUhyWcXlkCBfUTB5Wydy1dAUUi9ke
l5yOOK8NofE/2VEDrdveQUZH2IPDEl7Mwx883yxumrYh5NTvG0ALE47GYZvw4icb+pHUdH4EStqa
scdiaAJNfTf2HaawzRNJx7fiYo8lYBA5BswmlmEgjxZVMkSS/++8KNdUiwF/WnyzH+0EmTtZIMbz
8dGzYyQd/MNBRLlAxoZ9ivQRkQUlmyO0BraZZsGqUkKU6B6KQ1MmXZS29j/GZL28V6snK+KipHHe
fgZRx5wJ/jpdUXzxRYPs0oN36U4lGMLjS4iZfL/cb6NRGeNTrKCn8O3T5yUSY1QlxlD6S4Dv8pQw
sGvpU/qMX0NHi8EoRW+6Ad2jXOzhsTvC6OrQhFvaNxvdu9K5waqD9NVJ0TMNqs5UrLY0S8/eu0g2
vMNW0Spe3LHdf6bKN7qtlBTMkdyTVIDvxf0/bjYSuRq9xu0LOpJG0Uk3m+6tqwQlhgvZ7orfIJ0q
u0tNLom8vXM8wuf185Er3ri9fAKR7mCqTJuBX/GpOq79or6XFhYxAJQ77SlbVT5axNUu84jasUPG
GTXiVRy10MsBIAVTvar+/WsO8KeyhJ3a4pNYhtSAQe7xsQ8BM0NDAXFF9MQpBmgnL+q0/yhnJ5jN
+aymdHaWkS4FbV5mTKYXBnSmOWecQ6x4tEx4QejK/LS9WDlYGe2nWR5UHfp3kihrP4Ks7lG2YzLE
1YP2P3iHWlPpoJAy4G9MF1PBV3sE9w4mT1T4mqnQDg8/4Hs7vb9rX/Fn6tFsth/dIds/7xjOQwlK
RzFMbHMFwIrrzeD3jFQpMPCu3vfM53xyJu6vx4SgdPqr1x1X2AEISi3fdK3JlwZczF0Yz69lEEfb
wzqCv7rFXvHkvhOgN+bMm6oaX/lTuaNsNa5XM9BVzCnYV4/TwVuVSCUmnDgk6p5owkPBj5ooJhI6
TCjPa4VNeC36J98MX2yt0eSh0fX5yjUfxFKw8JBiOvU6alsY1uxKnrSN2q+rr2NSNXGOuaK57wyk
YB+7iJjZ1GkwrLLZ7s2Ff7hk9ffblcmGHiEOTg4/joqmUxuGkWGgD258cd7AJtxeC5cPlXqOdQT0
dRSTkt6nFk33ENm6FjwdzIJaiSiTeHcCzBzRzrpF+jMg9zBFC3lJkFHWdvq1d2OoL6JAehX5cwGE
xCLb/IruWFDBzivdoMZqRo/tbn/qJncQ723O9WTHBh6uznIceFKO5wSLnpqHw2EnKrU4mxTbbf9F
c8ITvhZ/f6xHczTktkTJIQ5FsFt7hK+TPUNWUEAvP2/t6gQN4KVGtfI0hz6bZVC7+D5gkEaF6cQ/
67CwlhPkOw5gBr9lcmeSWQzcK4J+BFKlhTmrCRble0EkXip9oV6B/HapM6Fn06JL05PhGFmvPpTt
dhu/Nj7O47DUf2DJbN+Xein1YHgYNXlYDXgDv7lJo4n0bp9JsRHNXESllsszRQjNJL3EePq0eEL7
cw1/7X8tCeqyYMnCUGGFue0y4FmBS5H4XzJj4PLhW9NE//cIyfQb3H1xoG7AvQ53YVxqe5XPv7OU
bPRW3lb0C4zyL5oSX28KjcgePQXBo17j0lCra5PcXRlncgX/fGiFuqn89yB9oZajruDETBL/gTiz
w0V9bL8As2zV+KFfK3L9NhDRNV8MsOzmjRYDJT8/6yv9RtktWSugQ97I19B7uPXDjaGahk2H85zH
H0QptTY2WSMYxBceSyiO3eA72M0OOxRoT05z7vMlcBlfDayFgQ6oFgF+EELO4ev27O9OAYm56qVV
KllZ6I9AwHn3suxRCl1WEHP2ZcH33BP80AOO+REioVA4KLJQDQSvODK1sbgxMIqHLL2ec9d6GeVz
1UaOXvdMoS6ZAYVVVy8j0QHkIJMVv3VqpZ1tu/7D0eNYPuF7lsvcSohh4PTCUbeI55WeLj7W085k
xlsfuI4DR22zthug7aq9vVT/KavlPacpfX0gdgUZUpZmndhjmTyl6uR/tFXsjgVO80Oq2Msa41IN
Jv+XLjyd0uCF6QQxD53mRV3JteZh7BuTG3BHjawFN4bxsVXOz3Jv4o1/RdBglKd8HGSyAg4g+Ffd
Ub2xfICYLwPIk2dKYNsyjNGkdKQPqzkaCmWFATNAC9atUWUtIYbYP823UNWZZZn/jfEbFfKNIFKV
+MZrUaGWQ+EzfQuOSVPzCtwCloviplM/phTBliKga7kWqPbE/9dn2C9E3Jh3d4WHoSeGqeeAZbqR
QfVHkTQMhguFzSJChdZcUXIGRttDN9kwtWpf7hpb00iWAFbDNbBFgwpSdFFZXeQtrVM1US0ZVCiv
hJZSZc9mLoGRpdQZ06L5+KojljUJawYni4mPl374dyI9EAySF1dCkFp+KSPlRs5vWIV9LKmduwsU
EPTnd50M+I98mPSAoS6LD2OJrhnOkcZTy1m4VOJFpjtTIeETecdw7LqDjuYvYYwHSdnk1WeStmBa
E/Qdsbn1f+8MTqcF2xEMsdVWroieGuz3RqAKamoTRSie2zjSDYVaI7+O/NrKJ/qTeRk2Xx4/y1ZL
3LZYu5x0RzvAwNJop+1kYRhddQND9P7ujI6lbGQk9dCJvbY++64bXMyXsJgiCxzQRu0NkMoEkprg
PXuYMwBFeB3AuWY0RtlyTzBnX8no6AseQMBiBOJldSicTiT2awJADn5IWHnRhRKR6ID1slyAjupP
fOzkWRgsrQoGsY0eQ5MZqnig8UsP+geKJTqnsM8vBcoEHMmMPMtxfkmWF3HaU22bjLAfQpA5CgPT
lilssAzihfJdgJWCsk2cG6Tqs9rdCBcLnIx1q+uiYOBFDiMDXiC9WZSdZKjo87DN8VtOXQvuYWg4
AwsvVx5mXOpy+rkRkEOD3MC7csykwbkNt2Yl4wc1wQBeoD1FYqaLmzkj9/2Av0J1LYUaCFXo983L
5ysmqJY5a/RiNybtIhhOLCd6hd381SwpED+gu+tF0W59F7bfKg6P/V7mvnEhBImOqFJtVL74J/Zx
eBM3jEwLSdUj5yPjAxRHw24R2e8p4k0hKDFo2l6pbHI7Q+iom1K6VzLIdgKdVjExhnpQmuO6oKyc
4H2Dfu8j1t0QVH/HTaAj2ZoVIqqGCYrSryIfRidoAbpPxdZKiZVum5d1UysLHm/erPpA5HuQkumj
Cw9b1tMysl4/L7iMiCpFE3er4QSJmbORRp7lw2IH+X4ug7Ecb4jww5D05r7cojLZgyPuOkPdeMTo
PMD+7OWH7/TMdIj19utDMPo58dDKwQj5MZu2uSM10j/YoNdPTFKlMvxk8wZ6BldZ53/VVEj7shbF
aNAfi4Li3pzW1lbcQEFFw6sz/YrZm3BhsLHUAXSA34bzoJYWvnXjvavWo0HIUcS22Vo/Xauyg+Me
crmAwcsfTpg1WINxVvqDt6FcpB7dB4qfE+aLZu7VS8r32/N41i5bwmdxq/UmxrTZKdKkjjfVMwfo
mPLlHxH3iNeMPGyw1p5dn0itICgwwGWEW3KhsYTMWOc3kbT+ROuLLwe5iI1fp2hbhwDP3nigB7XH
pMkFMhvZMo44+553K4a9UabMMIOYhsNuENmljSGmkiTxuA2AMjb7C3TAnvIFtguR8kXsr5IJBdVQ
Q/aJENrEj0E+N/I4/W0KupcHeUPkgX3iiwh+8lj/qzASPcI3m13vJ6woVztvo1Fd47xinuG207Ej
0qUxRGrZmQ54iwdx6+ZjzHCHWnxaMoBCnHrdM+pycwdBnCqy2rHxieDWp46I2GgAy4T4crVaYDLo
mBHw6WKqqdyZwN5v/63V4N9fFx+tmOrrLjASdLBrSHiH8VQxbUCNQmaV70fLNZxc+QWKsK9GxPhx
P7CBZyXPvtRtcsQ9Sx05wzx02Ol6ehpOmD+n4oVnGzGAwF7CnLIpNwg46od91wsXiOJtOKmtSkIg
imyxqNNe7Rp3CYsViIE3AKMIRoAWD0Ah9Fwsp/FfViV0CB8PCBgsAOvQvQGP1K+1j10sHfZQXHuQ
ss8bFnf3KikTxQa1x8ud5YpikheRhXCJuQuCbiW8lqbpZ3f4eHVvGVVtKy6jHbRhg7GxlizsoQO0
5b1r7gFvSCrnWDxvd9w2JDh1OQV+2Jqzh90sulBh0lWgwTmmCK8ksQfOwRLIjXFu4DgwIcV3xNBe
MvzS17FZ/Z836cET98gRJn/qXXXLP6LhYtixYaqpdA4Fg6qETSC+MY8Di5532bdcVaKd1VFNGhE5
36mcu0tSdpYIPIgBNcy7MJUfRTvyhQ7FJgSJBC1uq9p8fy8RZ0OK9hCdnQpHw6AlukWpD0EUjak2
H4dcGgL7Qp5uN1A7oNEPnjaWp+z4NPjYpBlBXLf0gF3DAtHxR0LNdKVAIgGGPNSf4X+Mg+/7ntgp
3/bHCQHl/ciikkF/dISCIcsvl3S1hvpz2aiXXNyA+LnEE8DIKIEVl+D2nVXblhEVARWYV4dKCJoz
l0X/kkq33zxaYwbYvz8KS9ZAwLgM+E82/Nat5DxQ4owlDkBAz/e7ljK8YK+Q/nIx0+5p1F8V+CXL
uEu3Dz2NRbb7yKrOEsU2Z9p5cgXW2bouKzgUF4bxKxdqVAJT5Vh6zrteujLS5PUpEHSmwteJtgqf
gBPcmarpHdJbOdUCP5MQ9QHAoCl+dTG0ijVq26NjnQ1rRr2UltM/SfXNURnEYLy414vGRJT3dBnB
U/CQ8FqAA5HY7xgyBp+dYTsUwGjjNPGOjXVFe5lJGO+2TbsjFxXD2/47vK24VlpGCpL4giSOadIW
u8LJAAZ941WAK65msvXCFSa75w2pSnYoWOfDzgfqa+CN8bmM5mHe4zZhw4Rvu52RY6mQ9yKrI1dj
r2itfJXYObtw1nzB0iZEbKNhs9eHmEazxgqXCB9Y7vNMITvtkQ+Jhv1JWRr5ROfg4Vvl05BckWhN
LTGPBYf/QkmnkbWzZ1qPlDWJhW6IqfpwkihidvVRUh4e+G/CfWI1Dxa5UhFDpT9dzljqc7Cqn+VU
dga6NLNEnmUHkKW1a5VpyhIIfttZNnxbjdxYYA3NgjV7frx8I9jvpxVJSZe3b1eT9XMgc/VNpGPb
TKu5DIgrLVpHFanyafkz6SygGqXtEK0Du3co9i5W2LoUZfmHRPrakBnLYXCZ5WwqI888D1p6iqLp
sVkrYTqWsVDeSF/4CSfgi1pfMwM0V5m2RcNW2MEM1nZxczlbWSsYHPL2PyfBxPZYdCDEeiUIZEhH
lXve24D6agjn47sWXlvYkuTwbqw+lT3QHM5RXk7VFJ6e8tZo1rbq/31WNMPZu0GubyllUYq9Y7jg
5DFL1qyfORvegdliaZRq3fBQzxcQbvvk4Lfr79qHOdBX9SBJ5Br66NkK+06G7CXJNEx3nlz07CYg
rvxlAuAl+En+mdydCcv1N9ekqN2K93zwKBHxWkbzrUPpeqJj3vLCZu2jsGe2+WOVhN3PL7vFA/xV
l7w3Jr+rrz2sa1rrypQat3MmXGnGp9Wp9fVXjfurlX53556o8mnfnfZyMNXw6wL9UU0noMSt/jWD
bCwT1bElTysYfx4Q8keFX5PpX0BkuH+o205+VyFZgE3VbO2Z5aQomvwfNQpawKEkEuEOnR+VW1ve
fpFh06YMOA/gJBIehVPTiSt+9h50S9KezMFZu3HFiPzOsJnAwMmFTRgcIUjGvn0ITexmgA9sbZr0
p6FnIfHitoWD6SoZYHqDIJd6H1HFNq7YCJvAN+dh4CY9tz9XR0AGaG4q/hbLCA60HHEjOe8D5kYI
IYdXf/L7abGf8obIIg2KZcJqKITanp1AA9tUadgQflYdr3/qE2BeMSFgYgmLR+D9y5eWcie9rZkm
yJPTfjxR2wV6xYpxdoG6p69AdYV8/AHsi+KjiCUblXzAt3qVRojoimrmGh1geyDojGPYWLTegZEG
/UFukzn8dKBjc4rcKi8+WSVn0MYqmLkV9UFqEoVTVL6yzjZjo9vOwEusv9C2IyFHuSpReHfZMV57
+IOwdx8sUlBsdTTQ7NHXHnPJhRty8uX9rGOJCxqXu5A7j5CoSKiw2tN15QlbbKZFyru4D8btMQyw
hKT09TqbmIcU+/WBsEFo5E3V+z5L1mwPAgJekH58tBSTubXVqZHY9tm9x52Oht0183WjLGIQ84rQ
WhITNMUzG6RobHtzwADI0rYRsZh3XcMy4/DRoSuaayE+M87B2SQpMEk43A9cpdOy7NVRYWF2IpiS
18wT8JgvmmWIQ57CiTDfAgfUe8g9tlEx0PTYO5rZj8XzWLZcp9LTXNdhQOoExTwanYtaVY/lzCm5
a7U87mCmB5NYfxCg6WdP/GFDOTHwMhBGxqMG/RFkM5P8Nu3GoeuKVBqT6gkWO9F3Qwdtiff/s1pa
32IpWcxu9tfR8wYtBY100HlqvHR+PjgIXhPKBn5BcrLrvzehKknpXSvEeZgIRkmmIr0oyJEysPQD
cgWomWHGbreirKhh0vqyBzEF7IPrgRSTKl7qnzv6EczfumRGMS2oCBKzLKwTMtea5MKNVrw91Kki
wocnd/wGVbLfvHVxafzyzSmJbfsn32AZgImUiUFSN0yPDBt2Nc4ApP1/88xZGmbVEku9kCi0RCDN
0jWZbyiCGpLV4gZPPNzXtRN9HDzd4tkyk/wfWfyBOQfEQboGZDaGH2BS0o0OxJ/IIx+SGmXWtps9
mpn4UgAbjWTjpD9gLAmJI2bHcBHbnA5L2OPFF85q3a6ZcjFqB/sPj3PTHbGwsPlpiF8yOR6hFGO7
9NcZRs7fgZlhfNPTt6R6r6ROiAggjEe9AZEZb5M4kWn07H1Met/P37NsJD56HC+BDDfekjWCiY8Q
biwNcJIzkgi+B28mbHpwWEtM8FzNanMTtMCgjbtqOvbB0aeXvDEQGrwnoC4f/G2cfqJqg99VjyJk
cf3JSc5Sd6UmAH65PqswocDZYel+UibRzNUREsbW2388GVXFpov1QTlwqQLF5Cl790ARo2sn+HN6
fR+r4wdfMwMJ82Wku49i8wUjMsE9e8LjZ5/YIP7+rGTzNbAtOGiHYHXd0H+SgPRP1aFs0cniQJNB
j3WZ0J48hsz2BwIYbAvzyiBft8O79OJrlHunZ/6nlBVRJRwLv+5T3KOZmurFy9bcRzWlgpQ5I50d
b1HdsaNFf1QFYhQJ6oCS8Xf/yi75HW0uI10SpeJCfjs6zuaa43HSfm7jiZgz/RWLCe91uar4jqKE
BVPmuecsLMg8fcQT+mDEPc9sMnG2jAzSFyrE7wvdrfp52LJDmaO4/yhD2P/pB6pF4XFRFN95eJOb
MqfgPyvxmpJ4oKZJWyLczRICvsWBspxPAMJrt4R/DhgoLgt6q80zj/Shvk6a9ifVoBkw2VKyx0k1
zVeDxy0WqIEsbEnEZyayAQJ70JVHQmEc9g7vCzLtaza0drk3KmrNxR/v+Ezk2gFPJYg6apAQbBaX
sAJdTfG3Fnfi3hWsAC99tRPNwReOr1zp7PIWozyGZHjuWwin1cEEJ/QvpnKF0GdE1g/8gpaAOmy4
2XDvc1db/iAlYGwLcsjmYw1C75FPDEVU4QRksej+4ND7gZxr+LzUp7BhuCpf66tTUare0dpZNafd
ZykH+N1K/SHMuIvY81Y7Bx+YbB2Ev6WijBMr0C1K8U50XA3GWlBRlCDwlk2tnMGB4oLqUXC40jaf
Mtu9dbbWoO1lNyYVnuunGjxcfFd+JS8TmgFw0zV5xqQdOh+sEobmVHnL/RkwuXfYqRnV3s38pv47
lndGX+sz4cnxWxPqK5+chSMCmYuqWdtDvY4sh4puu5W2lBOuS03rv6o4euV1hNFimSSC4+xGZwFK
PtGfWfUgi17RMKUOo2KbeHuSNJjggYIhAENF8tqVtaRvBsRPYch+gRUEXseOiDzix8Q34VeptPgm
CXHw7PDqyX3OXYNbMWO7/6GH3GFHmiWc8fkaICXeIp6rxnl1mkzW+eONXhGkoznag4Q0JQmqBRMe
5V7Mj5NNGu10WVE3a24YyVVZtoo2xk1FJ1aVfpa96GrcP7NhXBQjaDo0JTvHAyzrP1I0wi6m4Q6G
UTxooN9zdizReEzoM+q9qpSHmGYEFYMxXPw7pEauedGExfsiOmNUCWSsfBn9DXpG16c0dw+XvDBG
Aokk4y1cHkTJ+FHy8CVzU4RKs8PSqTc8pO/ERQjmVV9IT2JDDEpeq/j1zxnXKQ79DYXOnJJW7RHt
0jtdqqUoW209z2iOe0e5uSSFL17MObKH9CeLuqEa4q32zgw3CPxBfY9SN/E2F2ZalpU8HwqlNx8U
4Fe/+rR3h+VqMyqoHrFJMoiPHcqhaF2pOvGoQOxHpRMCfXkAcWDJPKd0hl895/o3AA4gwFUIrj/g
HctEV/CG9DAeIX3FVZ50j6ynJFGGRcWBvlc02OSVTeCvqxZi1bqHgSq0eF5OXOXp9noMQt9ffLSP
Y1+yZKKp9LX/WSM4h7qehc0q9+PHCohe+YEsKUk7CwutrWsJRGKyKmiAhrISE69agOX9mSiGLYU/
ZZw+WKANz1j260c7YkNLKeR4XYHxS4W7pI7EsMEPMKAR2/0k0iLGuONuLCVoSZxM+5SmucSu8Kak
7I1aoHaAU0Wk1slWmA/jJxbN0eo6JzcfCfXtDEoStRhtq7jou/3x7KMDuwAXh+N9ZsUPa4kmFk8B
ZtXWGVTLoRFeTrxwG2UqV7reMbwTbtO9TpYdnw2uExjXCv7pli7wHrTWB2wZgrpGGlOXIldkGeRm
cHzvLCzsW/BzUukPaH1geAojCX2/ntYblrQ3mSz8SL3IK4oTTudm/9PYy4X2zRmzLzGHZztbcQ9i
mlDZwpWT1LTWUGwUvESl7LclmuR2QXD7aNuaAJjNCJyJRdLELd0C9382H1T3vr+JPZSCzAghK0HU
z1RRop5UYt6fdVY4GUWKKynq6pJjvSg+0SP0C70StPhfTAH9d2d+vkBjBzL1cOfhBJXtzJrY+fO0
upcxFVrCWhoFnZLZR4pAIbIavVlo6tbvhG4dG3nNaoTROoM7k5G4CLWvyc95hNioEmniMrC+W1aM
GPpvLiWJg+IC3HKu1e7UtUDz2bvJHaEcZ9fDlz8oSNj+GW4DjTvcA82zrvQezItWojcSb3TLwCnM
09rNsH7XYASHZqo1k1eWi/szcu37vOrgB2Di698NvI3VOkWJZ2owaQpKdby+zmZWkrKWq6F2Qa5b
sQFuD9coyDjcN/lsgaB+x22Fi/T2PZoCtrKXXFtyd0UPui4qra3SMJSbv/xhSM7xeQ4J+SWXmMp2
D8r/7RrCFt96hXQRKZV0LSGabZn11fIpI5QB9OTLAQcTWnb437SnTD83TbqkAntEbwZy3uOBp0IU
rTMPuYylVFqNf0xzsoDcSuLq2N8g4BMOHQAhkC99oU8Ixz5NuO/Et6Xa0pqFgVCgZOaqEQz0oPCk
Wgho/Qk4YU+e0ixf4cFGWwKlZEXWwgJjbmesQbaBVKSSUbwsFdEDGuvAb178Nz8kSDBUkPq1JH2u
/VqrgBmW1Un0tdpECs9LpJps2pLenmcatiLQj2xACTe6FuscG7ktfaMTzgTDBV/cWRApZ83ooARM
QmH5y8MHHdPb5jq4r0PjsP2x/7S0+3OMYXTqDHKa5tMChGS6xYjbPXi2GlwSvRurVbBP6DwQk1dB
9dowB0aF+Qzpue7WEVQv0fBCoKCzZVj7WM2/9jAkHxlU662F2Be3QP9xxwmJSoREN+crW/Vi2JZc
1rLUdtZJAdRZ75Ka0QqqGXPOn9TvBPFjRW2JfvrPKXfyTtgDLWsoKgZxWaKxyYjdmev/x5bz1TUv
t8kxPg8jwoLblXJD3/UiZ9v0W45eUlv6V5r3MXXLBhAQ5DjSkLcCmsa55fwR4k/SXi3ZsCE8m2d0
xuwTQp0OF24bHhZ8jeCNxdUWqJ4iLfh2+VSdC92oL5Tyd7arSiGZ+Qwu8YbRmIsDhQ1F0FEdh52j
x2HUU36aHNU+7QUVA3qywpuPpT0BNwvgGCOGb6HuHZOwuL/1ki5IPVU2Wgp0HOrHqhdeJl2/x2pM
GrejOHs25Ys/qlDbWeYCCOtke/bNp/z/jLRVy7hahsSnXQHf3azlZDvkd/7ZfGmc8x2PaSsFHH0a
vxq8ejApoAf0MjXXEY/67WB6KPlo0JwNN4gywMhf8SBe4NbfbPc6RYhy58PUsCgfRZKY10DgKApx
/hauxsAlPedcxz+CuaJNmC3q3VbU/jjQAIkZl+MfBaEbtTDHsBciEzZXG5UjVkKUPayA3NtVVBa7
1gxcOK7bG6Qb2EhyDyW7DrjbCMZ/5q2EqwEaSJFvpjMBm4kn8vAOHjOSz3NFCn/IcIer8VLrSTFs
xSa7iX/9oj5nTp+/QQBdCUT1bypDJsFcMX0Uv2z0CiZcO6tqW+FcXxPRV3E3BQCzlnvr5D66QQcs
QtLcd05TD1CxJiqKo3TBgUkxCXdvt/cvGPlXPS3b9b+x3UPPZVsYOWN0uXQzUETqCEm52UKcV/mj
7EyDWVLTEzxRb11Z4IGZdxz2+QZ0hDP0ww1R/bWA6TzvaGK3liappkfK3pY0EGpwLcmif0nf2BDF
BC5SRqKl08zmw1HIzT7GcHNSdgyBVCy6FleBuRI//+KbR47KWAOTz3f8s8Z2KOXWnYQxStOL1iD3
W7AR2BsWTFUkHAFiHNXREJnBck0ML5hE0L9hUCgNWj7z4dfW9CH9qmlFUGKQsNTVXPJszUISRfeF
I865EiHx34q4oFDA6dTYuCyPtoYNBCYyF83i85jHRsI6raJ3qTH7jKx/Gv0RxqNOLkXjqyAr/9BY
Pb5Cx1Gnn6Qx3uC6Pn96qBlF0QE0Wq/9Indn/c4vKCaXx9sF55dKt8LClHCn8YZGvxcva25jjpxa
ARqKuPPMh5c6v3opiFJq8pbIYkS0aNN3FMO6TbBgmJYdhFMPGB/k42+vZ6DVeBKhDgVEbxN1nKX8
6E+33bMi4ZMt6hdOhE6LUjQZXYvOSNTLGAgRrAYkVgFmaKA/m1tQCX9rRxKzA9FRBwASG9mFN12k
nB1CtvO83Cs6JE/e76+MuA/dCA8c0XjPQxOWiCNQJsRSnc+8WN9tBP7CMkFgGJZTuPxJUYuz6gDB
VtgHorJiLK4cllGCp0bvdHjoGQq8+J/V3+0b3spzBii/EV/ZiUTyLulPibZfB1o8g6DrHGbYXm79
SuQOSSAz9shLf8W7ET0qccaaGlDTtd1LnW/GDHYJfhcps18RiZgw4hwU9l6g+CMMcp36nl3rHlrD
3raqqi/eJiUurBiWPK4Woj45Ta9evRGwHF6KRvMb6LqJQKGFP9wDJ6j9aZoa3b5lc8XVCzI6FHkz
2s+UQ91fHfGXgZCBmyHYLuxnsvVBTaiAjjJm+BqvctHal19vzSkxWelqFpwok/aKMQ6+NNpJTAbD
jApV04Bi1fdw1R3SrEO14tCzLunSzrF1M9/RO6zamBRUe3W5vqOfkW7G1Bx+CRDYp9uFUdJPbP9W
ZJDZ5ryondbT/v76fU3UAou1TzU/hrKNaBkBkqudRkGcYYEcWaimwWvqSEb/OOxRrmS+jcEfQlRg
WwXC0AXt/DVvXc4AY+Nu9dBYU0wxGqvUnYr5bkKYi7mzGDspx7ahhoR5EvvAAAhnwC0ST3WIjbOB
SUX3tCiifN91XJcsvJFNLyf/LNhK0Fv562WccTtmcl24kToTj14HcO5W017AHn6Qsq+Bf+FyDGF6
MKcEp3Fz6uXas7R1AnJi8JZQrI9WCw8FLyeJGCJvY7jsYVuPVPJWZocZlNrGfFktEUgXYv5V2Go6
ziOajvTTv0VjqHNhVWxEgTjoYj95K9lcrJtK8tdFqqRN5twCBgeclTcwJ+3jpslk2UML4IGg0Cfo
/XsWCxK1jYQK/rFuW2TmJupdJ5M43wvVIMAxUtG9+NCexbmjKyD0u666PyORkQyJdDBYR+fNwZgn
nIpM9iuEbLR+lBQV8HOOVN1JF99MIe8ZxDhW2ikspMNWhdurd3kE0hQZMDGSPPM9LNifzxgfH+8j
P17buYTnc+bAXfX1Ao6/XwG26E8lx6ftGFpAZZc5rY7k6UnuVrBGlU9GlKKvLP3d3i1d27sYv0YW
d4W+p3zZoPrs4rCu/4Hge4ytp38S7pRk2ll3AjpSQaXyu0axwdqsWZoMqs6LORQ6BoeOIqULV4WS
b+aVkdSr7KoyzuSfWLKgdeyiVs+kP9Q2MvCGhZgQLJU2S0Ur5RpKHotQlLpdcFUTKcaup1q3zylE
KKPkU140meHpf9emeDFqyYMwYqWdg827sLxeto/9ezRvW5NztABOSY56XvjjOtnXOUSD7DIvr0hD
y36Xnh8GKAOgF+EcmI4DuZ9CCUaFog3WxsjWzXtVtHmfJPS/TuNZbc7G2Wcif6wnssNsqvDg3HmS
m79h66MNXpQJ1Tre8USfU6zIIwRmdAeG6eN31hWFF//gch/bLpelyXzcgkYtqmCXf6cpwGrvwnt2
wH0T5bz2nSGpQlTP5Qw82H7DeRjG/1IrLDSSKJP4QmvpUorIGeO5efGDLDeOSJjMA3ktqoO1OTen
i+f8tt0pwhvXZFX2rfz69mo1LQP6EJJTQVXJzLbzEcRYjQOjASPtdL1RvfRH3UA/AusMRGoJMphg
+47ZFZqeDRkuVFYR0pOhhuUBQeyK6GKMuIWnN7n3iACShG3e6b+Vb74wJJ1E4S8lsXR8e8TcRi+g
JhdON3WkU0qD4mA+QmyMmIPO5qrpB6qB6enVFfhIhbTDTKfcj985Q+9TO4DxZxdvgylx8jYkTdsF
OBdmfiHs+4frA7BZouZgY534oERPZLKJZ9mM2/ADTAgYmYQKf5GdQDQRx662+tV+t3PNDyl+3D/N
C997aHKQZCeZ/0rzp3rC0Ifbs6z8Z0NNcvM6x39wiQ3OE+I2iAUnQYygOF4gzMKcx3ILYh74P137
LidjPlft7GDxf4y9FRpMqUEWYRm6mLVQT0RTss1Yve0NtWo7mT1ROLgQDv/I02ToUw33/ezIsHBy
PECJGwpd53yX659ll5Pxaf92gRhFkJT07lNPWt9WQIFwM69wkiEAf+sMweOy9dskjYzEU7toO02p
nKqIt6tkUUlWVYX+H+LI0X86v5LecPJ1W7zh1+hlSLSv/jddwSa6UzmSCumiRh/I59jZ0diQSXcR
f1nD98OLWsvCeaE3e593AafhqUzW/ojvmeXNIasVqfu8mNkqXyfLIMnaGlz816UwrVFKhqSS+N+y
tUdjarjyPDxp4EhMkiRrNRCbxPIdq+CHdPtb3rHl6TKWUptU6YQZELeB2/s8eF3QkKKeXXOujtNx
FYZtfiHEGP45qJHsaa5bUiNHawFNlps8jJJY8aGtw9L0VMH6dFmH84znTA9r/13HE7SrEriq6JlT
YESuo3RhThZtcD1mdxG32AeWxCLQl6xdhwYhVqheEFv7XjZhNweX9PPDn6i/ZbwJbKX+zqAks14V
RFD3qqnGwxafDtNe6XjrCx1Y029NHYNzwx7O/nDqRFQ7W5eWHXcDjlIhXvVsVcbDMq5UoZS8tlg2
n6I7ViGE7vhxxpgOOy+7NK+OkWirRwdgvR8bLgXwkeHhZU5z2RV5nUiqi0FKTU4gHbmOlC1584nG
Rqa75jOn4VNbLGDzH0EW70HhnwFSFnXBQc/RZ/CUJlNr/Q6pAB1EzcwezUcr5FF+dx4gl8W2UILu
w9g7/bbR/c9/tbz0uPYzme0TTmpZJ29xWzr43ZtyMW45TufL7Sd6mTmlFK7u7OWYSyBESiDDZL4x
cYKDMwuxF9gkF/HSEJ0z6sfxJP7NvV2cmhqGX3rC7cG0LLPGSyxeYcUbXkNbaAeEf7GgtRDJBGCu
O3jnvUUwKEXmBjg3wiplxPubazEqgue4z3E/eG7DWuVoOh1L0Y1HYvi2XubNImpbF8AcHMpvgh6m
IWuYLroWtruwmewUXXgoMIuQ4/iLcStC5cekca+IpIU3RG4V8ymicQEA+jeHPVE8iZuBbFLcnq7q
Ws3TDu9E8QXzeW+NnHLlbF1HIUdVkuQ+79dNvAkGQrzTKtkHdSFl9wHcKgqkAyywOoVQ2s8ij0bs
oudopvqq1Ktb9kh+CTRltqnWzMEu3Wwqy0dIPpqkv1gA4yaWSKNJ+nyd908X3SPI3azABaIjoXVO
PyjpvMGDPdLG4Ss2CbQ/O9HEcj/Tn9DTdn84zgUGYl41xCtw7ysUamj8KkwU7oH9wcJrvGMmvWCX
Ct7F24WAlFbgdzbfyrEfLNJ+P2Zq5TG6vksveFT/mMV0F/4Xiq+BLMHkQtLn9ScUngwAG6jequIK
FUPZzL317kLqpYO2TfNUaPM0sZtGWEUW2O/IltNWQnMNCmdnSLTQO6eqIeJm6ZVepeGXOOw3Jyfv
OnISNuwl/UxfQDJPbspr5T1Zvo/ha3Eavol9eOtTPnwp4dJDuFFqUzAHrcxJUzAIBlZMIuAj8Luo
kBLRVZVdGU23VZv7+PYxOpoyFsaFa/iNvO6c9RW8qLSQbxHb0b0vk1nxzn0q/cp5zcHiV5P6m63r
8a4h3M7U8BwS7SXzplOeu9Y9aw/PZ51rXiikyPTLaii+/iOW95UAV67s/kvjjuabcvL2fr7zVKJQ
nuHS61s8EFW/Cq32nSlTgPN0dzmIfxbwHCBIlNBj2yhAv8J9za8RUckq6qvKuTIn9i8RTS3bvsuU
r4H1AWemD3oNWK58q9Ioe+t0aaPcpv4DUiYbuzLGpR4s7g/TNONdBEcNFooXdhWOkW8oFu+alEcQ
NBh7bOsGC3GhNmxYCyBxKLBIdlNQP01drKTHEkqlKbVwdiai5Ok+3Dv72yZJTymokjBPfaBD/vz8
db5WLhbBBxcZWgMmGfF2CJJYgR6elH1z/lD4SamLrrTYFoCagvoMsjhtB4SR+V08WULFXMFeqPMe
tBsLN2wSs6bNlh2Q9cSJi/7yrRgkIc5o+T4Y9ZhSkmqY/XEwjjbf7QJuoqePVnLq9CDpSKq1p+Ty
tEIJWea7aCXZebQxrMnBKKQEMCEHv/fRF0eRqtCOwk0Z+hjp7tszrxxC3o71fdgH6bwTXGjddhJY
hQ5uk8V0JxnKYHbBqLWMt5tiKp7sUJw9duoeqrSty9SgVgsqEXnpFCdcW9DsCFxz9Xod3+TM+owk
67J9Thkm33iaOk7whFs+hqMqM1sHC82wHaVuEJcut4i6jofzUP/hXZkUnn7MJO8GUDvhazeDT4GW
So+UVwDqloctWyk5waqoVsV+4d4LfsN8CHUhEOy+4wp3tYwr2cecwnEOxbGV+FjG73QNmVsalpHg
ZXNVcPClZb97YrtnVpnd8feC2FZ6dJMzz0stTgXrME7g2Yy90ib6VMK5i6Uuu4mowTGvZu0mP9fb
FCi/ulQc0QdUO06sQucaEjRCCf8UtfgisqHi48V7igepUsRYmVFhZKjWDVnV7TY6T2WslgXpmuMz
Q/2IOcB59XkRyHUtc8/QEsVxm9hg1Zd8JUirev/1g5Kr57IpZK/ioJgB2k9uXX7psgeCOFgDcXcx
UzUf+Pt0oDWuYRpXKZFFAhVKQELSjnNQqB8Jf12FscOrwPjl+AKeyRMpyS5rqhLE5fn4EgLFJ7Ms
q8bzHu135jF0OY//Dxl6O8pAsXvf6ysG/wvbrvLAISrPAJ1PInCOdJV8Dw30g89cSN+J3P77Rrsb
p3sWBf/8JMiyAERTkkItNE7JUIVhCAqYjDNVTM3ll8aHkzLr9vaawcN9J3qKL5P85N/WArT+uVyB
zxhTJ5jopwMxfHLJq2k1VKcm+zMJ3L2RZnLqGxZjT1kOBm23vzzhZzHTc16LRjvarGcNDM1Tcg+S
/wyg7BUjyvvkIYMQ03ln/Rv6gLNlIqRmjvVbKJ5OnUwdt6AmFwTLcs2KEzshqDWTrCnyJTOUlkCJ
T3oUStlWHBNJHafhEGHsfV2ec+6gc2VKjuVhceSYKiHqOXjDqjpraev099cgTC8MO99TjJnJSQsI
czGeuNdx3lQfbstHEkcjoIvpleHfNXovEh9HFWQ1T8LzQOEESuShaRFzszXpbHoWWqSHUS3RJt6a
RJ3FzkhTsXMspvD1wMHvEB9Kt3QzG5KrUokGR/PiFhWv6XilGyRY8CtDA1sFBJ3I4fIcGLM3dKFL
NrTJrtOBFTXQlWgNWuDxOPIbKPqirfqEWbnoABTdVXfHfaQpwP7X2ne18qqddv++S4Rr8PF1duId
p3VC+uKIkx9ewC+weicxU1GaZ+h0KrAHJsKLr/6IyW8JY/DrMFP3o3tshvJay/FqbPMUd0qQpFgx
jCDaFfyTz3Rvaci5T7fHPKRtjH00jD66mmrKkhFuErIVezTWN9MyUCn/XaDxzt0smVK8CsuQUKoa
yZF85vgsX3ljN4XFF/C2P+i14HpF5mPaEhoLg0q+IATsSPZwKklajUSccKhflAwhlcoCSy5oUis4
xr3D0B4KtP3ICIaXeJgTrYqDVAUjaXOa1vU248Bw/DG42sFtjWW3njvdtZNhPkMKn/ZrRJAsYrfw
xDAYWfcmkJfHCJVNhHVaS2MjmOuWAx+x7xlHuKDbF/xakB3G0Ukl9fDfsWjSxLx1krSCGjtVzUCy
h5mEcxenePFMRCc2+cF/rHUNreKDTYU3SHKRW7guU/Jz6etPfKDj6uu79IXr3wIcTXHB2PWtH2yo
YTrdZAooyOwgz1Eh4Vie/pG60ZMR9nZceiHFeCstiNSf4XSSchMxuSpk94OcWc1Un4AqXxPlNn6X
XIWL1YhJdPP0XE0vBfMBWre6LxcWX6j/TiBYd8OpHNOz3cOgHtIufC6Q4AgWx/w4x7/jltG7T2vb
S0cScwapvJU9lgDogczB5k/ze1kSNrj0966N5o+WIN7h7U/LjFXAdxo9KmyjE6M0RdYuy4vHXeqA
OrHZ+6sXa/KbcWRtNjdUzpwdOKDNkDcWEVWHH4BrA3Gipyu10ycmMXDN4eSfN7UNzMt3FNpu1/mV
CN9pXZ84GTN0Kd1h6ZCswnyZ9NBYIfcMAKSGBoXp9tTUIc38l7fKwYubbxGMTLRqJLNRDePOrEku
IifGkbaSXoxDy7vsXuPNjSJYW6aSwehkRqX34OIeacjgfNydRofGAivEKyRxPcUh/zvGAZTpVM7y
ZccxEXEZ+DK61tz4Dim08PoaJU6ftx+O26TkSUsiYLp6ytfzd4kRFKHJ8KoDk7GmA5Gvm96VVL73
KJx/+ov9TEvwnweF+QO0lnyLImJJK+JsYZRFJJLwxWm5DVfFcRdqHMfEida5GMP9ByMqxloEwmal
QNpK1FN2ESmV0cbVnXYkFF9TiXVRRTN0jbEM4DdkGQwHOiZUV9NAppwIrzXcppiU66T88dWyKn3Y
CkQHpQQpO1G9qBxAM+esHuphO3VfOHF7ZTbBiO7ucJZKbO7bJ4oRnSI2sPnqFZHGt5FqZF1fKcWl
LQm4hTfAG8jPU8lG79Rd7uAvB3/Rou7PI1WufqPmvGySlymStT1fl/JT+4SFDR1jBPXoJsjIUvFk
6QQUyeVXxaT9V+Dii9tG5bRPkMsd0ifGngEvJO7iXIgXEO/PT6ldZK7TvQnnLMbHbFJ+pLOctGa9
Lr8zZM47D8QTUoaf7MVgsyRgJYB43WzbTOnzSav5JRlhPuyfyBW5k/e5gGq5q1aUIsPH97DJ119b
M0rxJ1wAYU8CplEeYyqm45q1goNEdv2kp9KyBRQWdmORqf9gPgotK/Wik68w218lsYUp6L3KPOaD
zqHAKj76hqRT/M/7KrFyaQnxVUIV1dN6yKUA88KWkueua8PxnJKEn3Yb+FwoUL1mEikrRpqsRGyZ
+6USBd82ngg3JB1ibS4hNQUB3929ge/V789xaQcqGVOlIwCTrIFRIr99q8Cjo3KBJ2TFM/vrzdeb
FMjmZoOPIl1sGXyJCAFX6xFaMh7YwqqFZ0w4FHGDl3Oqdi7+KEsdYG2UdZlBGDebdFtM0w66VvrL
Qw2N06rF2BPA3wyI3ccSk4BZs8UcYdu7DsmE+h05NN8Ruiz60oazfs4o+021TLGRf/MwDM7RiIcv
J5R+97nDCsrBwfPfn0aXpQkBbQ3sY9G5UK7QkSw0KG4vAxxDFXWUAl9v0oymPJric6dqf7EtJibG
iEGm3SvJhqbiQgmPex+J0MUtZwIQQlyxrPG+P2mCQmz5/6oCUOT8Yj7AgXkOWtqbZEa/+NDzTWG4
cUXpmne+WJKSl42yQLhERbMLEoLdvc25zF/qio9MmEyGSm2oeaT/+rdcYCAOlUs2GNl/+LJbg+19
Kjz943eSjn7iyIqHlxMv65iDjzNN4QZq/KLnazwY1Z0/CVUkF5j2IqQHeQnaItN/AtJDQuCUoWbE
75hKUOFLcpBIF/hUrZz7COSYBIoqjCmBxY8gjWHMZn5Usv5UN9QF3etQbphD+39wAG5Ljs9z7gHY
kyQKUSUVh+W1m5TTJFvTZCqN5+VFZkDLkMlZiSELugsmt4Qr8SLYxgwUDUt6q/EC0L7tqSBiUJEr
EKw21zcPs8dnu42uLUHOk6gtAdkVUru6p0p+qVNnXcMCNPHNM2N+Efv05sGSODdTUKgmJNcNnO66
HqE10UIH6KV4rRtXO3o5QhXyV7j42EIkK2Hlwp1O0HkDn6zT+jGz6W8nlaI0Tv/pOUHJ6o9iNDbU
GB0/37B8bj6BGKiJ5wm1dPLnEFZimM4NnXkpOmPgx70jVIaMiWIUBW9eS6Dy8oeYWh/lRWt69eA5
wqQj7t8SCwjD3C533Taau0Z0NNqmW7d8ahqYHan8AQufZtWo3gFiDqo2VM50/8TmHz6DUPhEz3cS
f2/V07ic2vsFX/5AOLYLHf0HdgfYbBxfVWKPOw/FzzUSINAOCqrZ/jSD5PPTbG1agCk2UO8oQ/Q1
p2L5sgACi9BuuRkT5WW+tbJ/NIqK00UFHrnWVaw9zUfej669ZRx/HxTfZfqLJeaV+I51UTkTsMMU
/VaTbO3gYNMP96jMejLb5lVXa6EgUegx+XCv+yJf2QmVJWgS3VOdVSMXqIr/fEOTnZpHdPwXVkM6
HMMswcu11g1v/PrzcyBZme2yJ+YuK/DG80Vj9TcxHVLi4NF8e3vHo3ERNblJ87S466eX9gaifUwl
uQKIS277Y4Rj1HuL3lzaQQdTVGPOmPZ7HkK1IgNxeekOck1D8DzKVjWfnBoYadGCcR3A/eV/gUsd
HoNM2xNgJX6qx/E2gXuFVWaulLW9HJYf/DJFn9lXrElel1eirN+BlLgLIkddnzCTvg3w/sKMo8Nv
ctZ4tKzPRc9i7PITrfuY/DTmgxQROcMz2FzEum/F3hZO9eVwasixSW17SBK9cyse2jID1noImKbr
g9cTiiL5o+Trq66MEjbI1BE1c3Ou2N8X3K+d+h67UwRtB6dKOrIFffj/LA9C8RKKfP1no4F4QF7a
fTpIfppt+qcvDTSsefC71Z9GW0VFxIJzEmXICqOy63O2xlAnwko/XFhFHQmP63bGqU3o/LbsYkly
bB4GL3fU7hZTdyc7H7xuz5lyc6U9Wshrvg3i5mGoKRAi8b4U8tGD9AOfsDHyz43UzxTdIUrKtutr
Z/XuS4hWLKVfX+nEp9AMKt4rwByHLuDseiFyj+x6+OsbXRUlchIk63b4wU/nH3nSLs0hltCps3kK
lKzTwwvfFSijwpwar6Kby63y9IH5REOgD5eDCR5MKsT5XRVUshY2hD5iOXx9Zpqs2Us3q0pJ9z1b
OzzzHLvRRtZXuKqcbq4JfRUWiRjray1Qt7c9l5O+eB/sVfd84UkHOV5m60M9WelmbFBCeNMHre76
/mwte8BX5WCJTGx0XaSN7bByVSiMy/KCRZDj/vGK2wC3+snl2m/a4w9Jd3e+atC2rFxH6R8+WYu6
pyGScmvJYomsHxyrDk74ElpQz+O/9NHOFNq8GmA8egfj/mIqwJYEXOd1M4HhuJBcEqXZpj2fMcea
qZsuMonQgZl95rBcvN+hWpBhbFaiuchwpscsPXXEc2m7c1LJWOFTVie4/kGuCtynKr0zZq/g6yOz
LYlKLZQGzXsOYcjWUc+j4aupNQKeNshe3Xt54EiQ0cIp4qDx6CQ2b7+HPV3XAGtCB6W5RvCvsv5b
5b94auu63j5Y/DUJPtXgXDd3wP89krkkoiuDCbA4Q/FEyd/ltny4ML5nSSKAiOYH/2Gz+DOnIW0D
xCKJr2xdjhXLoQvsklP1jsq+d2eg8RSTPrk2+BAE/eEc5SiQVXN7on2OgQ28KYB42cJbkNVolZHE
pTwd9aJeenkw9wY53c5aqYIWTxtNWVx46HtJdchAAe9tae8YASDyfI3YAs10qz6wLq6r6sLAdBGN
EHmoUL4ohpVGZ/Y4HJV+6L3+jOajZLt3bmn4P65PagiRWmvtPXsqsUaV0QhwOFIP7kGv73UagDCA
F72MTQLzgNLRi7X0Go885J7boIO3MIhiivvgLtX0kzBizUREn6/yiX8O/8wciG/QJUx4gbZjHYI/
6X8Xc+ocVcIaiWBZve4LQYKdyBuVBHqoM9o/MNlJtYZJaSFvq74TrztiJuga01gGC39s1G5n/LSB
pVHBVOtePONpDese3yC4VW5RJuSTIJbkwgl8q/fpxXSEM4G4oxveg0MDcf5jpJAkmhThgW/NWFQo
jkgU0cfAwlRt6yGL7gxlstUSM/EkwidYkOQTBEy0aTdSVm2q+kUgumfEeWLtvVz7FaEmn5eALkUM
cXCQ67FQ8lseaeE4dp/ik8GGl/TQRy68WAJORYNH8oPEYYflz+3jX5tzrIdpkbI4CX96OGaOwaUl
i62P2m2jklzFT8B4j1RIX4yad8kL8s0fX816FHQ+uih81BOHAUqYJak8zZIrIYtSwAT1jx2Xi2ZG
PyXKEg3NLO2ki4GMDfcp68DCOdzWrKe7HWFwWmSduifgQ5sdLoi1WLfvycrWi0rukfTL9RHoMJ5C
FinL7zJD5+TJpcF4QSHxNt2np4YU2UzQ+kFfyVTpVkeUUppIp+zJzKhrjqaonnGemVLFV8LyInsy
FEKXgUU3Jk+NFA5gMUOplZDPvjGJXXeKUc7t13DE9uEsiKZfIthylGG5wtXUAqUP5DOkHmmNSl9a
gNByk6Bq+cCIEpqEo81JuEly6aRKV6zMam+KnUz+5Mc0tOxgRv+4rW5teVzYFvrtmh7MZDZyAscs
RV3hqEInctXITwZN+AdO/NPfI7GxhR7gJ1xMk4BL/tmD4V/lqn90pi6rqQEtSztd5veBFYtVBzUW
xIhNpkVvcq6lw3eirFJnMmoMADq79e6V8GQfEnX3Y1qs8cPHbsKdyU7N09397x3fbQbwsUyLIqn7
yIOSjO683aDzUYbB6cXwcsmi0u5oR0KnyoN6DPf7UK0PJXI6ZAa46qxBRF9j0KccaJL09MtFar7f
MKCbP1/3Q14SCGAeHDRMxNlppPqztJzaleuKYQp3LjGVCwF6YDqBP8+o8HXAMwQhNplyt0++0gab
c5KmLOOE7rehOW0or0EQGJK7tAGNNOPjohjknoTHd6wKR3hiQxeTozqtjvGqVkBBQFf5tPNtTiIE
Vd8R5W8gmn2tExlEncoFBg8fqLgLFzn/gjjX2rN3qsOn/VGha4aWu/i9X3cz+JDtSkeNOVT5PLon
+I1/Q0gpRq6d/OAJLRrujZx1XwsHIJ7Ie4Aadr4kEfcSKOftHLP11Tmk6Kud7lLJ8W7ndSj/gJKb
c+ueITudN72qSIkTMtuJHVtpF2JaY6+DMzhG4R1aK0ilhOxQDL8dBThqWOKNVqgxDC7RrPDqzs1F
pYqAmqPktgxUxH/YDw2UsQUpKf+wJChao+uuh0ZxKPOfy9Uf6vNa2BCV/n1dSEpIpVwnf1f8++j1
Jrm2GqbHuI6LvmAsCaBwSmvzA9sU6OozXn8/dBZTMmjeEpqR+GoRx8oSPFZGcQ+kL0FB+kIZQ73u
1rluLmI5XQ8YqdnCRjzbz6lV38XrCtfLaj2M1oFF+ttOYrPmtj/ZqanGs/yN5aL5R4u9M6ezkXHq
PcGlbyK2ZrCttBZBa/wTZ+TNrbO9cBj348yHPQ55VykfpTTkOfUwRIqICkngmBus2lkfdTUZ+aBI
T8N4UuGCpuob/2i4Lp0U4gCoBntDnh9KYbBDWw5QOPe1+MmhrP3fbaAnJVe5K00JsB7YWzXL49BF
ye6e89lT7mR4KlClzd5TkKgBGcZR4CUt5Nu7jIh3QXs8N3jNj4naXdR4Ck7CY6itM92kGzIyIoz7
FjZtsGHTc833lHd2/AOZCdxo26NzGgJMhBVZzUPpN4gPIwOpfn3i1NdFwOgcbuBIH3hJMqX80dDl
qyf3T8mL4CR2ft51HPnSy9QdG9R45wJooIAaCiL0jSmtCegho26P4CbHiuNvD51zxs/85pqWwR4i
XHY5UhZFa8MJNSQBXvFeyuEyTzkW8cM5Emzxv3q1Qs7/sj0f3I/kQbIaeR5kUM31x91/I7MBhbVk
ktlGxAmptU5CgLYToT1pMJBgGwnsEUCJau8qNu/UoYbHc2xSH90gfrY0hSzSroc8n2vOBFftJRdi
8RoXqfnHaNEJ7HJVndGk/B5BgZIGi3Z4/aWC5TgjOaxxbToLt4sWt+CciAOx5D/dsRN7dgYjltks
xTc/bq7EF4C7/Sc02fjTX5fkGD3qWkiFWCMfihSYYM8KS2Cq9EZuXKDRDhNQ3qZFCqNoZJOLV8Iw
eK49eoojkwWbyON6NuexLAK90jmXzXDSg53cRmO2SnMa1h9r1rlJ1sKheSFQgspr2WSOeMDKZr4f
K6h5IoHZlzMcDCHz+AVKiizKoTqEK7O7yTK6yWKbmT760KjX3kGyUcc9zG+/BwGZQ4KZ03kXKSXp
Eoaq2PHW2I4jbIc35gxzTmFF+JVeN2YSZ0+GrZT8yOTWxNe5ca+ueDd5eNoLdoYxPaLZmiTfYD0G
Owl/u0yjTcweChSl4rLWvmoGWBYTeAdJ0HTfPqP2o9m2V70FnDfquJtiwsccO//bHxLFYtpH4NjO
UI/gtD6Yq64vrr8ajxglzSvUiw4nqxu+qyE7li1hKtIJ8PmUG52vKz4ddYzjwgQSvh0QViN72Sln
4KYqgfpTd1YJVMVujC8JIX/HUQbpG/MfuhR0nG985qvpc2KFyvysBwSh/rfhzaXhN4cAlrHybWdm
9u4zu6q7cDuHbqmQau5/E1wVgeZQ9zO8X+pk4YuiQitzOvFRD8O/WQfy31yJrIBCuT23AcrxsqYZ
2gLKjqbJydhQH2giof5DEmp9keE+vdr9QkFOe7InHyvDEbzcmn3ANn3RrVL0dvpr4+VwTPNL+ENj
g7AAatkkY3MFXREwnRX3et99kkVSgWe7dKuMqI+fUhccBeNdP0Gbc+bVgXRWw+W8cSB3rN4hIa/z
T8etfj7Jkwz5fwi5MoxU73A3xo5WgaLaxXL8Y1AO5GMCuPk+/VAPEb5/tqIba1sURDxcRA3sKcuu
lTcIkgGYFkMpd5BQe6sMDCnvjZaYX9xUlPytfSYp46XTpt2i8rgA4TpxLbMtwbkZTTXPK9TLnpcb
HsH+4wdhU0J92/kalb7fcIs/L8BdWH/u7ImJqpS8CoqGOzSRYBsOoKALH2xELN/jWBCjd0SYNFbx
Rauc4wpx7YsCJKOKT+VDz/lodU/iVrCnscGGNvrAPwqy+CUCUFdDIo+2y48T+bigOOWXaFvwnjZH
4pvMQ0d6Nr56oGEn0V13T3bNbWYT9wGa1JGeJQh01p6YdRIc7t6G93CNBVO0a7jEQyYBK7gipEOz
gKEqOb/XO+m6dzgah2Ro1IGjc+P0N+LjZyCzmugc1WRjtJgsC5+4wKHwtoQ1x/y56eOiEMnG/s6d
C7Nueq9vgbeG7nnm0BqOBAIE8mebRqdja4YiFg5j3xz8pN+DkC1M4Jb4nNmYPTy4o/bGmpQc1D3+
cNvKQdbHuoziaz29c3HA4oQ9a8XWtsS7Eqob3aEadjxWI7Bv80HztdTZZt6nGws9XTV4r7/iTk0p
fqHR7SY17wHYuD6J6RNQNH+NZk6Nzl1i6ps0f8XffGif2CV8/iZEO0u1wYCnPSMQFOoEJ5ONtQ1H
uC/gH1aw0LNn8k9HZRcNzVCJ9NI6fjuM284QSJ1quNnDE4J/HXD71pFt4MERiHx2Ehi0G1Fp412H
+GRSK/GNiy9fM59tehnQ73tIBd0DyPWSukWGG2L7OwSY22ZX/pLTGjnalnbbWmGVj6inx0OGf2Zo
qYCbUPRuWMle1XP+rC2D0YedqHIMczCb0hrUzA1KsbIc/ETt3ZJaDbPFTsmw/wiCW55/D6/s6O1L
4zFI1itZTXYCux2saxYCBNsluT5TJ+bb6f27xIvD8/N1Vfiwsq6REe4RP1URyrjCbO2xHeGekwmO
Cx9TYnmpmosZDcqy9OOueNQpm5XUpGsAvaiMS6z4+C23E1mtTrNda16u67w4bAx9FS+g+c687SqT
otJ/987agq3gNEPR/ot76u08rJG9icpViA9hvqPH8BahY4ZvIjA0C2C7UytMgqRo4ji5WydGfN0g
nZeqHd7YCqO4gUg75XU9lzhOlGaW799Y/uyzueZ1oV4p6x96BeR+IiF5YEXBU8NNJCs6sZNy3zFT
p6K2nO7/74prCpaiI88DZC8TtWE/zCovSD2curOBBW4PoqAoerxIrCfpHnU6bRF2iWNiW1dEsIIG
sAuiyid3+nfwtJigID7k+3rqq4091ke5v2ZR0mBHUQu3J4eoqImCkuojc3S2VVRYOkDTptCjOppz
v/S4RwLNqoXKzn0i9CbADO4Xd4J3eUO/nGwVI0JYo0Tm8sRI7UOMrYIw/voDRqIGEhSJz9xf5arg
Hfnn+AJT+6IQtuv/MLZLjbLd2OK5WibGCLKDiDa9RASHAC58ZSV3JY3DFlFY8U7B8t8HVOOaTF3e
lIQ6mjX1F+Ow1bRsfgNM9eufJYrrMSP7xASqUZEg3gOcw3H+xuoFfI/+GFF8bZM+SLiesST/xirk
R07TnzLAOOl3rvAJndsFxgnvYLZ+onzeBMcDIqgqTI7gcPap/gr34WxNQzcCiwftV1jZfMGYqrvN
XcyyUc1hu07f1U74XuQ9DaViBx4AXzzLzGrvfvUOkz8DKQc1MwnLbi8OV3WuZP/9gvEN5Ze203S8
MLfQ/5qK4rYR3a3EvpXStJlMP1sBrB7YubvdBWQEi+XDRfnTGYcbkxSWT+zwXYh/3XKTe0TGt3Xm
UGD5DUIIueEx3SEOhg6cAtzZT/oMWUAVFDfQ2JUylSfx2CfJJak9bV9n70vp3WqRq/UNQL4KHpPs
23AE1NIFORADSL85dJ70Xij/nurb8sT0fZK58qarN9rIl7pkElPQmgPBQXHAylNQYm8nzLhsFWyd
C/dxsI71IbQvGhC5IEpfffWeMR8Srrt+dtfY3P9Y2OMyHV3JcUQO4sFEc4meEmWdp5KNoiAKdvd+
bjxXcTcejZrWt7TTxZZmoCskq6swW+c91Upc+Q6zoB3xsWUbNM32ou2qrcJW0c0//j/cm7G1ozGa
WHK+CXPrM3e/VtXmAaNdzLqy3tK7FXTVZvem1h/OhMS+ECIMf3N307qDpdEo1pT4w/es1rhVkkXn
t+xt42ioQutmlQBPAqj9gGJPiciPyv6Gv0QzyJ3s/eaFgqIRxrFdJUpkaqKmDYdYgUYvqwsXpHq7
6e0wDsH+bnp2DPiR8mr9sxt9wk1qNoT6pl/UYSrd5UDvx90UvTEG+iJkUPvdFTdOmhNZaWlzz0C4
uGn4LLe+1B3n6akQrjz7BS7Qxe/i5/C3f2r0j0MxhyHbGTvAcirtdRkR7VeWDzEdx3AHuoBL16Dj
tAVFa4ENvEeCzy376dNHagmXMqi4Ao8mY/KBt8hgoZZOVqEW3bcGtbBsZOfRdUQWKyy+642zg3lU
XbZuYwqsP1FrLVi8Gwht1gLcHhhljfjJgwW2LhXPGFjGrSu+YMeEDEN7GgBohdyupzI5oYdx+vtG
ioeAhZaTzwAP0taRyc3WHzySvD7kwve2L+2+eE8WaKOX3n+DI6wglAWvtzkaZRTN24XG7r9q5btW
bIz/LnhZ+uFBJM+FBflOVZMXc5H2d5+Hx5YfVpqBhuXXHPaQO8+d2uaKBPzZ9K16sqqL261iMtM2
tTCRpPp68kocku+n1XXu2I5jo3d9YxFJrxKGDRRuVXiIoAPLOeOjIgwSv31KL0IsQubaHNlxuC6p
UaVPIWz1gxGkDGMH+3p4hEFSUXYY+f6AYG4OZZVr2dEqX+mIEbGrjcNyNG5q/ZJlU4dC8tr7q8Jy
0gMNHnr+T8rVhf1WCVMW042VCPwQDjfqP81U95hpIs8Pd7lCt/+BXBurkenLgxEsKLvZr1oicFeK
LYAUpqQ23y00HGkShupHL6aIMrTnNLTg0ZLV2C56rnOSlKBa3b62KXCJ+8erV69L09dp/iEpkOQS
YpB3+e7ZLEVD9haXowuQzK7IreOIa7n7ecPnhAB6Pi+gI84YPbyQztICTueswpj8dVsW347QMoDi
EhwUS20jNfpU+SCcCJK4m0UUHedM8C95KdIqz60YRQ3G7aF5gM0BvzPzcWTtegzhpJQMO2gsfB9S
AKphK7UUmO21/d+c9YNdcTr61rBWJx28uid1fSmZXyGZlyJi4N+ZIONY97bMabqMWb/E4tiHIrGg
YCqaPGaq0D5/TuvwDcEylb2dYyANpI5OklrxDRV4ikkGbx9NevtnaNB0/XnCONc8SZ1puMBYp+ls
ukAmKwSKuhCn0YD7lF4+OIucdmK1O6egx6jydgjTjiKDKQqxWvG3leCI9RJjjICcfXLqzwGf3gnR
1ndZkx3JEv+pfF21A+o8O8z5I/hl++nYk7REW2rT02OmTHduGKTtUZtgjg85acX9T59ejbyrhIAq
W9ziDjwe9RfybkUei6ItoXRZR+l8hD+ZmwvDNfn54ikrnoJgQeEtB8HTWr5c4czg8qrFLHKiY7Zq
AEqW7beAdS/hBKu8Owk36XlOc/Ibx8uKsLFtZa+PXoM6WZXzFi+LM8lFB1QGb/NiD2+1td4iNuke
9oy8thRqlUo6Ho141AsIZMpRl2GFDDfGk8fvT6mXVaHSFWVsL54LVKH52sCUYEYFI6saT+0JfZJj
1vuOYJF4EAkzzx4yvkMzR+1gNbnQNe/cl/xPbqSSRPLeSaReiGAm7+2MLGOQyYpn4cVMKJdG5lvx
iEXQ/Y7hLi+5piuvCNUv15KsMfRXtSeoWZs4KBGFbJqBE+jJAxzluP0VM2+BwFuy1tR2yyS5LCDS
i3UHO62TIqtIIbdk3rg0W1kTGB/uzuHJdoUes+GCD2O4f3fSI+fvF1dHKmAJeJAtk8+FY16I1Vby
JC7gcSaLPH1ZjH2ZDZTtaXwb4id5L28xDhH7oUYlOyGlQeaAFq3QTxCRN2EOzSAjTp3OuXd7LTqK
nw+eO2T0cP5I2RLHoY4yKfQ2gMH62PtNURnXF+si9UNm8gxrd1awFV8YpZOR2DGDItcYYAunXfHF
tZtjnvTI6tDJNjTWoTJsLYXvEe6OM4dz2iG7JtfIT3M6kcgRnQy9JH6BsGGzglPcsEsEBDTpVk5o
RNY4Ad9agbSuK3QpXhPOi7CmLnYaQC2x4++2U1ZNONvjRyy8ZRfyz1loNrO072djVlkwHHt88jrf
6dDxVHs2SRwXyp+2g2s25qsz5ikBZduDVBJYCCrxbeX5vhvXZx4xPs0/lTuUR79ekkPoJJy/rcjg
F6+EzZ4dDBU5e3FxiL+EgQfJsx+ULW4xE9Q82dwjP1yM+IT5XX1LUvPYh+m9CnNgr1e1xUE5rk/9
a8mutjleXo+STqIHCM9JAx1v+WgUqLGoj+ON8Ph8L9BkWsyxiWvcoGkBmqRGd4TlKUx85alZ3UBx
Uw7qhzAgvKRZ/UnR3aHDwQnmKj5FVMLLiJSP6V4lY/LrItrSYkdfzLJUYk4v+GctCsNjijwpWdp4
AJnMQEk/QDJivMmDvUzpsGSCLBgEU8Nq0P5F92AQEjF879zBT4Z/22eY6OJmp3Uw1lmhYtotZ03k
VRCNsXZsZ/vQC+06Ay9TcfMmAwZzIJzPR1XUTAcfmkSm7UwS/QfO4iLADb41j1u19wuiFQqcAXUj
bh3KuhyS4tWhEmq1vZCtR1elL+SYE1nhrA/iUNKBfjhgAICLbK/QMG30maheWsyNY+KTWeOgFJfj
gBwsHZAAdOYefjkp8ore2mIK11DscNJ37geOnNuc4rcAxmThiucdMXUkkMb2jWj8yqCnCtOhAcC4
gMPVwpL4LhQr9BJTviqV9ZheBo07foaqH4EfqJdPd+4DcUJyvnOT2EbaIvhLNenjKIJN+pVG9g6/
voPKkFzGtCvcQjm/mpOvHKkpiaDkxu8n1Los0ojT1OMlz00R/1b4aNpLhayiSWv18I7ZhTNEaMVC
9NvsRZJPgMbdehKjCwFF9L2I4kKgB9wM4FA5XE6dgcRqglFnJF+9CsI6xEJEdF+kBYp54GXnl7Db
wCGyFkPTUy9KsYgp6e1uRlBKdeTbRUtqI136B5N/yOeulYNboy2F38xA9QLBNdbJsm9wJjEp3kz/
Dwvb30c9r3GcGOm+n9E2GSL5EFUiYEZMpZd5wVwF3kFCNtxKusY49eA3H+cAKMYSgK+SC9e/hY1m
Hs9FL4x42NvGK/LD40UeWxXdDUQboYu8WuWFWmE8ZEj1MF1PzqyH6J98vDdJYWXr5nj/5S8UCkIv
3VadrGBqAYzOGTDXsgO0aas/kAzyD6+UtnFLdkkDmhPXIGZ2vJkND4lYU0PsCUzZwSxv4UMuor1t
Z5E1QLMgValjdzbrtYNUeSP7z+XUBad0uDyl4ZoHayD8VMEEej4ZUp6bGIrFbLS8O6PkzwhvE9oL
jCcW179FcocgCaC5M1v2CP9H+ZG7n8NsK9Lc8XY04ZU7KGRI6IL9tWrHEgatI2oeDLxYd4I6Q8Jl
Lt2eYlv8+KbpUA1OPrIilpMLH+cPo5L0NSHPqY0ZKUMMg8c941xoYdHdiJKYL6ssN7N5jJXILt1/
HWHQ21qayjNDrWDv92bfAUuMFf8sd70BrBOmHMiQudeTb3Ie020E6DYTaY7DWZ+uEMVMLv6EqqrG
3b+ZwS3PYqwxqWVcXwiSzkfVbiqwxNz8izR3jdEXF2nmus4zfWGEWcgOQb2i2cM2V0heVTRv+gr0
jcEQ68El4+f6vRlDuf8Gq1tOOMJFF/ARd+AoVzUkEmIZB9qCwP72vaiJ5rSunx2wYqtT9edY4bOQ
8CcLH0UWKxC/xGkAS5pXeE2br+36vcefOE4bPzgiVGvnCIfBE4VUYmgIOZwlBf4VotL1PaHYgGZ2
Upp8c3kLhEet7DL5ASb2ZiiKVnMMC8S1XvNUI6x+u02cMK/4vBn1+JGT+s81gvucUEtJN1ixkThX
CP/gcfq9d/luDNBMnCM0u/xa7yMyKvJTvXx5Cep5EvFDgGEVraeX1E8RMCR6EXsrPUZbWbuVumMf
GO7jO14JlTyz3K+2FV6Lrwmi9zH3yANolYHVlLV883pyK8ca/NkSaBINdxhy3LmrHe05zHBqUIMU
ky2mzMo7wo+L0uijITAlMNX1/8ZQPDLRC5jTQFgyzA8y1hFyCpvt0C03Ci1tYgpNGhLCdxWh/abC
Nnet2PvEuzkXhOQPiCP2T70TcWtx6EzCWByFQo467exfsw3XnlaMZN8+z5wCZBeni7bpxbNkmH0H
7JKU/vQQuxtAqk7qrk5Vii/hfERns3d8bIuB9cg5gRgNt9KvO9eIDhUkmrf3mXfdt0F5nR1eqPZA
5SRpERldzE15yPWYUeFYJnJC9Zy5mey6vrS9T8y6XsxSzUcxtW+xFfM6flHI5smtFio6JB1qKO40
5Np4nQNhAGU1rlljPFxsmL7gyeVKiq+prN1F2Yx4eGRQM0yCcydOMYxD4hDmTQU/t80THv5N41Uj
OfJZMj+8ngHzbqB4+k42udULkVkfIvRtDUoqQoWNZdt/SPiRJNsRFMlLtyUF6AA/000wPPkFBrUF
iHbo56nDyjB1iDl7C+4eYVl4vI7bB7t7X8r2uJASUH+HJ6DIchD2H0wLhprfpp+4vD0M3nQFQH06
Oa/ItwiWgXomIW0kY1ZuYG0Wp86IgMCQyEEjS+qV1GMJhRy0YP6U8uVS2n/7xExWtK7oInVdFqIW
vm7JJig0gYJDJf1VcheM4kFa92v375zxtm/L/y4+8haQgzLzP0J1/ZLkYSUzxJeoYm0DAB1rMb4k
2ze2sATFITb0rtrFrf2wo7ULwMw6/0ha1KFSRM0rDxBWACw9nwIjNhZiaP6rC5hx5w9AsVOnt2RG
pbVLlYg3f66vUgPxg988Tp+MTLTv91OsTtcmnOERR286R5Z1NVJrD1JM1fI/tNnns1yFXwR6dKN0
PXBqvOW/ZA0/OlVpqDz0jdpa5gSgbfF+5pJ/A27ucDcIXp0mGaYAhUuemlTYCyQwiyOqWy+6a1Dd
PDkkzJQ+F73dARqryXsQBC9wUZH6sxBYEeC6xPMddUagdPn1Fdzju0puvjs7Xd74W3R07fP5AdkL
mgazmnlIDg1R9OXpRR3XwAA5KuMqvHNsIIrV5gHymGHY1uou5s1gV2XoRgXs/PeTUACSmwtGf1BL
P2R8eCINOKKmhPrH3EA3EIm6Jg5p5uDX6vECIM+bKXlC5STCh/xBKqrJ63FIV/SHhmbL7S5Jvx7N
52E4oMXc5O86NzakErEyL+jKUS6obHDhgaM0kFhotF9rVn1bNxxYZvYK/xavZPbVH4HZ5LnZuB2J
S9D4VyR7ZCgmOhflLSgnsEA7noMxFv3tvjwLbt4ZWyx8I6UJeA5mab9kTn7thCYSAiPP4Pwl/4IF
PkMcIPyWe7sn+TyBZhfK08uvjTvDLuf7OZQ5cHFZtKxTMozmc75HndTQ7VE4MQ5yOKcHyPuIQDB7
p7atEsSzqOdjuShXjB9Sq9xgs7vAakUt/uf9D2imQ7d1afiHqX+7A/KMJ/QWKFwcD6YWa/FuTZmM
akSnDKRCRLfxZpvnkIdGv1Chk6Rrl9Gs/3VnS7JVh5KEIwQGGweLQKvNmmVSQhPv9bERrvmuUHNQ
F5Y40+KhS8IwiNNjUDE9VuyLZerWGCk4QwO32urUKk9htTvYSVSHuS+AVJFqN1kmKeT9t/avYibz
97PaTE7n3elwhBuxvScCnEU6WxFdiGNoFlFbV6qv6Ewrfo7snwjEwt7ASY5MRW+8kAcLvW7k4PL4
xFZ5DdX2R5iG/T1Qf/jdZAjNGQRk9UzzX8NVtybpk/s1Lo7wnMjYNZGWpIpsVzLfSoD9piNlCTSr
FtAYWBNfTtZg5UCk4q7XgJ1Ysl+LqPFiZi6W177V6reg5Vmj3p6TJzAckfkcZ2rO6N74RheuY+gF
Mgk/yPvoHw4XoP0B1nwvID4sPEQidxws9RmrKZvKBRDdJuF4wRj00Ya4Dz6Gt1WgWHhq5dmTQLRb
t1vOMRx37NFr/8LC3aGN+OfF9e2ONPxEaDAMHgN+Qz5WQyQkium7rCmPvDoTa6MpUSzQ7I6xblFO
DaqXU6xQ6j8OGy4ZYd6UAqe7wbi+3UsXou4iddH+Gi6YT/WJszaMquoclLuKQSFUQYcyNSElHNRs
SVJ93vXIuY+0hWCPOGl3uhfuxdxDe0shX8eLl75ARh7FDtAy3w6U3IJyL+F0Rkpvbel1c3/DStF5
6hVZCj9pihN1gocghcHZSWjRd5yU/a69W9YZ693jR3+46xedfjOivCsUSFLzEF2qIrD1YLHaJVzf
4uGwRNaa3LkS3MBnzmpbrQIQfdhM1dMhOEMOvI+6eOmpEBtOiTIfc42cMaTtfJ4NC2OZ15W5T6tY
b+cHptPyH7uh+osI6nwFTV8RBcF9Vnj/xctSZSIVHUI+JQ+7NKTyh1YtaRTwkoybNABsxAUnLHPC
+3h8kiU0aE0qEd/Uz5SZGYay0mmNj84N4bYOC3D1GOhnF1PZ68goojuum6WJ0zQ1HtuFY3KL8GZc
Wir4j3Vlh/2Ugo0Ft5iXLsw5N/1EThvq8fIVXTO9XEEntb9eHnIr0ZXZGfGMrJeBijaxNIvzu9oV
RU77ZIEmO2FE2NJe5A+9TKBMlri/nJCpDbUySKzvuovQ5djA2MJ7w2goyO86/2Kc3+hPPoC52Pcf
mt65kmSz+E3U/agN5NeUevGhIhVzwhnVO1tThFN0fzhktKXZeLOwzyWh9f0RxNyL3jIB7coD1uBe
WYz8fe1U6ijVyGZP7/B+WkGIGflAIJGgbleNKIZHAZf+TQ5V34FudhmmZiiKlqqTcSGeifbtm3EH
1NomCnQNqsW8arD3iF5CIQWiDnaNTRhVvXKQfLqFs+8ZSRzc+ENWM1S5ctWusi0KIOb7QaYXHPEj
NxmEtFS8XVf3xHQaI4vBGbRi0KGmEEBHtNG+51ZN0uRZMbunnr456KPg3pv209difuudqmWlml+p
OSWh4Dw7KpITiGp9qNaZmaQBkcJo9Cb4hJ685vnM9k4NI2Z966aN25urO0s1NoeQAOwrKJxJ/Us9
7uqagTJ9+u1VVrUbWCHvZRGNpTIyAFtSUrJR53bVwTsV0ttEJAbcJD6ItWPB4N+gKs1ny/sGtZzQ
G7FKRJeZlFOdM+B6Ai+8jHGdou2iFqYAD08Q9siAvRJvQzZ83nIMkdHU2DSez86PGo+tzJcwFvYe
Ocmncq1foivMQ/ekRBx7h4EX3dfz5xboEdWnIRwp2jOBTEtZSkftyZKYaX6fxePnFExhxbwZySQF
V+zkBxEUPBsPhHlLcYVmKK2kO0ciEotBq5xTRen+GILu2wlkwDLup/3RtTy0kJhRYTjM48TaeZ/3
9uWphfM92p+AanFsql+9YXXnArANHECxabOo22YT2nVmpQLCmbvqDdAEZ1UVsG6iEl79GSAhQHqy
8O3f0Eacj6XFwE5/f8DavtX7sWlV6Vnzg5DWcqiYbbUuj4hEkWH4+FxExBHIwa3u+7ygFdFO6+OS
ueiFNWsnqR35S0v327vxZDqxAycuP2xC6cR/B8iM73ev9D0TovbcvalNazUGbVkfKg9bFyhbSpeF
dG/utEzGaTviHQnuOduHUwdYnmgbPUN5vAV4WMrSprwuYEmK4bQoPXz0Qgynv8qjupIjp5tArTeU
dWRulg5bQ3UMfJbOsfYQpZJiSkbCFEVbQKWB75ySPyefbZR8uh/N9j3Ew6YlSJTWbL0bfoPsQ9cg
CwM7bu2vvyraGjc07r9VLhYsmIktPM/1kxTJv0OnRF7mVHB1VnXI4tRtq+gnR9f5mcnsoWr16lUA
2A3ZocQCEDCuXjRfXPvVGz5QRlSuwjxao1kTuf2aXoHtkgDZ62T3C45s4GK4GWQ7ACoBv0VKpNI0
nRbXtlMovXX9NWDbANI4osyy1+B1npx9FIbck/ZMhi+VfqfDX2IlrizrGYJ0jjICwimarDpXP7oi
IBozoVknfIbS8a5OgJdVPqOJ7N7E41E3ksXX3FKtg6niRacJZzZsQmdlQq7sg/oLmFCoqXhw2UNE
4vaJA3Zez1L6g+d7sojW1Hw40kcOnsNoDslKN7IAWK3EVUFt3gE7MrnCHifrynYrzmH3BYnDvWs1
ErkwF3DjpYUkHHBKobARNpoloUgdMG4Lz674K3uGw8/JrY3uHF8b2sueTF6z8Tgyhh8sRwASq8Vg
I9UMnU1MNgQDy4SL2vzhKuw+5bSm4AMznbTY0na1cOq+Ahha3feF97rptTF8rUkkAGkNos6OqJWy
KeE7Onsxx0ZOJ+dVi7Adx243imUmBAPUT5KehdX9734MT0iF70JMsUo8LxJbFHrxRB8sQGExpOEx
9kiZq8OtMuH6IzI7fef74JU2GdLVoeBKq7Xvu64C8xW4AG+dUHNivLa2W7/e4wDiIoOqQvv/SOvx
9YoaL1mvQnZSGEljOAeuULD/b2VPtDsI6fjxt2C0fqKgJjTQcVOoF4znVGjaKeexjQTPLQqSEIS5
zrFkxp9yO7yuTD8et31dPa6lp7ZANsWLGOOD7DgKBpmWZKwTpH7wou+60PPs3AUpKfj7gluLI6VY
4DwXYyJ1hBF6jGfuOeHAQ2eAws5vcun0bvWQXfjzIcTjBu3MxPwDJWvL0iAnO6CgijLtaQsGq+tL
Mt5wvhfUMCtFpgYkDyT/tx+Le7KGCg0wuS28eMJiaAhgGsGnZolg1TGBi6E4zZlTFgrUTOy6Kfks
f6ENit537RIdoo9bc6KzbWJr33FtB3brrkY97+S9x8xfA3BgfaiMJsUdt/PUW92ef32ATdTkGetv
qkHj+VeLV8kIXXUGBuPml+KcFAFzDBPOE78PKmgvcTyoEJ+FRNM4r+Pl8fJz+b5YP2hi9PwQI4uk
CY2MYjght0Lhm/3eF5I6e2ezPrXkKWKkI+E4LllZPpZ5p2ZiQXmRkXpGO+duBCDJ6diDKrvzBaiX
ErmhfRMeuA89iFNkqHu1gwjHwcuDScMKBpIbrul/jzqpu3xT/yDJk13Jtun4w+7R6TighaJLlkZM
0dISuQQN7RfLSaveN8bv82p+mCb98lVWD/9V3NN4/8ZtHCxCi4mjtIlzs0FsHEInTEb5vCbEPaBZ
CykZUMjmqyHT4Y6xF8IM0zyUk4ohvfdPMgBkbGcroNNHGJ+WMIO4KfOdzx0kED/YNjgFJimTOoDG
3vQtg6B0+9vz7ixbQ1Rj6I6P+lk9pHZegHI5G83kgHhdShtPo8DyFxMMluE7TeEf01L3pPDrlwG8
MBVDo+exwR+nAdKBpiNN7lS2grHR8c+qDjNNxWMsr+W0F0AfCZNoRci0hVIpcdGl/Q3+ly7mdgmC
YYcAErLQsuC8fPPRUzCmUyyTiawlepB13Y/itkWtWi5u8/cQOsYVyaVNv0AbCTh5CGMamD6RnWjt
zabQxkSEOYBNKqt0UFYYeS5uUEYNSRrgG5u879TubiWJzxqr+I4P5fvWVaOvRYj9LaEW5SM5erWQ
9MONs3YiYiFKMhba82/vI5HAxIVTOlJrkl1+HHwJ0w4Giu8GXKZvCVcALtJJiaqWAkTB+QbRgRUx
HMbNFLVHy+Ckt6Cus1DZGnDvL4pFsqufIsLt/kKv4yzYCErvd9oAkLnXk4rma0shS9dwL50RaJOY
YER/iUXKB0ndx4DbPhsrnvQjtzaC7sTFq/lVI2HG7wJFrV2m9gfpyfiYUj8C/F/4hMf/caJdBnAB
KH0kjzPEkL1P+uN/50z/K2XSyAz9HQEN4qhpCOm0YXQ5VXcdc7Yvgl1UbXFhbc1RtXF8zw0Uwrwm
2q/dCO6lFezERVKaKpJVRIzLLTt1b3C/vZ4C8vr5sYJG2jzPqzcKuhXpjl4BQDDSv+/LPaBL8znY
JO9fWxE4D62JOr24xEwfR3yeMf+l2R0AaSzgPlDup7zF3UD5fFb4G2tJHHluEf8r5RCbWUqutG2e
vHV/jOjg3+/XqKToS3KcrMcOrmTlUveOI6MO7+GANmT/cmzNcVYC5MTezonD6IbXHejAOqXVtOa2
U+KGuxHsazkz/YfOC3U0CK8ep6/6XKTvRvmH9HjaqoepOl/bXmKX1vPqw+VrrM2gylykMBr8nNwJ
AT2zKuz49Qoxh2AosIYOtLVLSd3+845STqO2UhA8iTLHiJ5CLtKHGAbiWpdLch0fK8yugrwyQR9M
xSEZTxKvoF04lLAVvhLmanNfKC9leqGoI+1jTHFTPEo9MrZCqT7UHhzA1IdkJs6E9EoICfGhlRx7
0eUgDU5N943tfIjyg7S9knQBTTv2paVNJynS8qTDXd6aX/9gov8GQ6jsjWOrVaJ+ewKaQU7E+7p9
popGN3cyiC1OTdgiBQhS10W09mBVki3Kc2Jywr3ZH1NEj4/GVsrelXZVeZ0GOyiDZ//ySXJIK98G
yBR3lYNAMYEbV5VfdPH73mWSVtOVn4NhaM4907Z2xiRxEdv0yb6z+O7GioAG8SZazmIfrfL5kv8D
PdwDddFVHP4FekVa8kPMjcnHJV668Bs/qj81knKn7TrYYy4sop+DuQ1WKttazTRfCRHZluWgmit+
ImoCFQFUInQdFfhZBHZsfn1KsyLbovwNAzGQhdw0ZrCYBK8Rg3MmQFeTvRMzbDTGr1aUGOBeij7F
K4fe2W3Afp5sN/ubEwmi97XtnAFRNgKw8FDc/Scc5PV8btrfPasN8otm+Jei3pq+kJcQC+BeDZQa
F5YHJfEdLSSjE0YiOXzfALvXNKvbOq4rcNoYbMzuB/02QN+IbqL3SYGBO3W0TNWjKoGIIQuAn+DM
tiWFDmN+8qDRk4pALoJanuFf7fguIYlXkwMnXJXuZDo/LMJxif/9j2Uqr6M5AIoyk2yehC9jOyj3
oBg9IyW/Yef8gOO0RI9Q0P4dj1LgXDoRE0OjQktdB7CFcXO9ON+5W2it81xhyI02asdPEH7qLdzr
ODE3y4DUcJhhkUCQ803nr+rBGE+nTs0FUZhj/bP4fUeZ2T5bIs5sxwkTfOJG+GU3TBwD38xsaipk
e+adUfJqNKKsHhoOuLiglw/mcGx+rtMLGLQguaxo2QaH6w+GvDsIUv+KJIK5kydgxAz5jJ5nfOcd
7GhfJcgyWVGis+VJ14xF88xDwrlPcRUQJ9KCz8WiztHEqwo1zN255LZUaRthpbTe9s9nqBJrCTZU
/Mq+rhQU69o2wGeDpu8api/inWEab6AZAY1fqXDMea6sN/UkVJfeO/Gawk8IsGf0vvL6/ZhbmOA7
mk1BdVS2e4maT5s0MKAW/Ft170BMrppdc66gWmn+1wVTS4XoZLY2mPxHSVIdGIu09R+aZkZW8psD
IoKH36LWDUlNe4/4K/sg02Q/qbz0ZeIR6oJ0Mq8OSdYxSVoswzkDdmdJ1jQPNN4r0AKrgzCgmS58
TpU8BAGG3dYlZ3E0Er5/qP/GoaC+071wc1X8goznAw3DMiQa/ARmnz6/sc6+jEFzTbbRJEQBZMzT
NADRMFJe8k3J8NOjXwwlOke6WSpryFrKdpRIlwA85yeH4OC6Qcyy02RhszzKaaANPgigu56tujWT
TZqSBIWhY2iFSVlN3DYl/lTSSxie1U6ztELsZ1MZA0+tNxwhK2UPxZZTXM+g8KfRjo2jEveGOTE3
8i7FGDl3senRaW7awLbB8FLut+aLTs2nHhINd54ea6BX3CXDRQaGXyaAgT4YSMBjBQCJ48aqrF5F
lNPhQPDJ7ZvfwoQ78jb/otZJDc23HoS4kE28Ttcn6Eh+dLGHfUfrGgw8GgiENqOgsKLQn01+BmUp
O0R8gQ3sMlA27lJQGCBKiNT52kym1o1HoCvKZwJB3C2DuxgZZSueuF3txG3gXOJ73/ev+6PjlXm1
DWQtVRlmwAEztf856lYJfLCStzi2mp/w/D54Y9TdNmtCXBP6TEbO4uRX0CZvEzH6B3/Np23hVwq4
89aWbr9+s0Fp0Iu2yhMIOxE7r2oq3VSpPCQR3ZZEUhceDp1ryDOdIpWheOEZcNOQmpHTphP2zkKY
zMZI5hY+6mtLZpWBHan6hnEk+9LRRV96znknEnA/n5xdeB9NLB6EFHLc56EbCK6IWN6f4lYSdjpw
bWMUmSHZmkyaR8wxGl1j/+cn2Xqr07V4SPdAu0nSKWtd8qDu8LyqjQsbYxiyKZ6hFarf0O4L3Yxi
rMIdH2Jw1kyJdbebz8J20XTpD4zbfyBaoFH9AGHk23i6JFbGDsa/FBRkiF32LeQSAyvuV+eRlP1o
wn1tM+WMmjECD5TTQXm8VO48EdU3h/KWtLe6iqM54rUDKwpODS6l4lyjdaWXPmB85iTyyYhNholm
NGbn8cvA5uO8jWpaStPBTZMzucz+qlw8wWUjijUbFAnt25qNL7lbXlBFZohXWmwwbmSVh76LIEhH
bj6uNIZ4YtOOL5hLlTe+JC2v4ygtISIJwH5Q/DiJwly6C1I0QQaycBiIw+lJCT3w6GMpZdcTGvAO
0BSlFKwSuQ8QGsHGFjsDUt5K9ZlrmowNKYJM8YIx9qmBfMAxAcoUpa/JwOqz7Mze/DnKcpsyPvB7
jaBj5WkW3mZMdfrHdmmAshbDP84oSiK1IGmE3N/4TUdbt2aQEgfWf9hci0ufZ5BWAgspyBdfkhhg
17VlwkMo97opxAFFq74hMzte9rSiJa1BxrCJhoohx6bscYGlDuACebeeYpVNN+jKaJ4JkKCsrdJv
QUsodPyt9B6ITrHpXFy56bklYexwaK4zf1tnrzoaXBmahoeGcfO93wCxvlYXMUK0ytc29b290u/4
9+YVKfTZLA3hEV32uiCUIkFTb/RCLCdsQzLt3zleRGQE9AmUGU/PqASpnJYwmPXGm1sYG4YyzvTd
umKziGX35upBjefKMCgxUMniiDyrseBQ8KjNlwIdSVvxqhs/DVsUAwlDNkHnWDsv8v7rpUtDgMnG
ygA28+jvOqrA9eH2s1/wnywM1YEUX/AegnTmFCtTvaZGN+TVcJeorHh2IrkmrQ2pg/nB+K2kGm80
3SGocVd4ipqdv/NiKNk28sEPhE0iGs0dkZHqtk646w2ORG4GIpRw2LFceFDdW5RFVnX5MyAWEjQz
4ENWMUPVD8KkL6nC2gt5gG4vOM2OV6YWx/1Us9K8ymaLgQQSMin6zgdaAQqj6doufjEafyd2s1dB
/p/UptosobOH3Q1XW2LOKU+ZZYd/ECLMWErAabnpS+psLavW8SBuEeNGIlkf5Z3I9YZe8JcpLQ13
N8n701C/hRROse8t0rkSUHYhJ56g0xsqt3LuXShnNZkPY2yroJjoXG5gAOdJlrt3RKjGCthCZzBo
Jw14eggJev3D0Nlyar8T5wi1DtKo+SGXBBDpA7bS002Sz8WFCYR4eas7Kf8bjmnLbcmp5qu1EHrV
4nOR9q01Gy/keysgsDIp2mHH4aZfQUIh5wCTPt6Pb+C6qYCrUtWBHoVnpFZTZyMguG+0KMfVyheD
aG71wYcm7Ih+/Fjd26eQLo+FzIG6d4pdZNplF97fP/u9vkPDGF3A+ZrfSUHcdYdSxP0yiQGubg9V
vbqcgZ0RQqcFABQOiYb3zcSaElnnOLC7oBXitsFXXS38Biyu+4xnJKRD8B4d5dLqQ7AnWejDutto
AG/H4v/+sYIkiuU9Lfk4oCFb31h97oEfbsgo+0GECvKuyTeiJ3V9DP+PsLJdXbgdSXHWxvEf8KSi
7/4qjCGGxE+iH+rLotEZ0lXi5hY9WQ4WuSOn1JqcCwYYHJOjLQSwVi282fHjnp3qFd6RpzUmGCar
wVv4RikF+hUmaauJVMQ2UM+mlNMta3E7Jedf6ussAkswZeo4AiK8IbSA6ZAhwBT1MT0PQnsYXsQc
in3SeZTQQx2yP5Ir43hgn3RPJ8dqNd3ZdJ1QCPdI3v1pvSfBiZeagJwaHgs5YCe7UqbyX2I17UP4
Znq/c2d09RYMWRuYQXv0U2dtbmdUHVcvaQLVW1IUdhxL0erylaqlo8ZjF24sU5cQ1+f0xD4Mq68d
D8arMgn1sDLp2lecdLFaEUGsQafKQO5k3iu+l+rfVkHBYudfKHqMdGaOB0U3E3bZY+MJ/jzBHL7g
fSc24muF38YROlQghXX5OUUWKC94mx4qRMhxiFUAJzMday5FcVC8+ryfGS/sKnmsGlf1wF0CeRis
wdv+9swiPkicXrqGkC4rd9+D6hoxBKMmw+9wwxvAdTloiCjDiqlPzuXVwc2PN6IEORVNFlEsCWIx
oyvRHFH9J4pTAKAgsn69JQTgwnlR9MxxTkuERuM/b9qFAEK5cf88wGcaEBeeLtURfuh4tYd7t/oo
n1+BU/mEVbYaem07XwGTa59YA/5Dr8tVinRAaD6ZpumI2AiPpXVc/XyOD0oTzfvE75JESG4kCgsm
kX3pyGiGT1duKou/EWljHlKpwhqbHmIEvzd3EhERB7suXMxiTyKAKjPEIbOoY9VJY5jLj6N+ok0g
bx6SEbtF5QXoVu4jPPcvh4VjgOqBnd3ao2k5oUnRuevT/GhEiNhifFgjogOTLMjLGNTIWQA3WgnW
zUyQHnBLPT9c+XQYJNkMZAU37dk+kdajrK7IzZ8l/yuSpZdT/q3TRqgDfcl4pcXMnbd9BZquuMki
t20XNLAAlpPHREPcmcQkomNWqtsEo02P13JnkQXyRux1j7QGpr+Q0AitVsDoh1PQN+9rLls5MnbN
qA7Wv/DKvKL2UMOf4uvsVfWtjIBbAEgXfvgNUHV9FRS6XARJ2EcqkuxX9GCCa+pyLwfbNmK2LvFn
Hgr/ZTRVWshEHZnQXY1Z4Bkms28MaL3N8nGTwqGEPU2utGKk+zkL1RX0sHxRYsNW39roVBvZPnpx
Fh4MjvWRppRV8voo1b4Ty1UXV8WFC+GvT2rGn472Y22dAtNX5wXvRVjw6fmRxRYoMWufwXe/J6jn
9RS42SWj6f/eHLF/kCzKft1NqY7m4YpkMpxEjRb0itY14GpPxz9h+nIpUO7I4MxSgX3KYqD+Jfko
FnggrXIeFAxBfe1R+jMxGpaMamqyctRQxIdcEiqY6l+XkWdNFWKS3MykX/R0j7tk8tVg0YDM4Sf0
2163Hu5Hmvjk4N84y89wQwIwW7fEHEw3GB8qmJYIvqzJpMpRbKzsktWEeXtbwQueALbYzgDu/iwU
A0az6tgUwZ/Zj2fSXLZT9EGaJvTP+s/zyyqJFmEBZqi6qWdBzpYmIObLR2x41YF74BqUcP5QNSv0
h9tXqcsjPqz9K0o9xA1aG2R891CH/sn5J3Fom9YpQENrG2w9lJx44FYMAjKjk9OtgtYRWRWf69XC
fAwRkJ2T4ytyBipaO1UVpGhbzuWn7+W14RzJyglLOa/qOfQTqeABvPPqpVqGBC+PPwQDQBXjm4Eo
4xxgqHrjZhrurDWURSavpKVCUM8YFWv7312iyhn2RLkquwM/lJ7qmSLHrVyDWWadUS0MQeKONM2E
RdeZRVgOUyVWp17BmrK4gRkJHKpSS4Ys+cxf0K4rx2DOIlc2LKsed55IJKwW+VFq2Z7+80iyLUs1
KTQGQWCLgJpan1ORDMq+J8PiMUm9ruIwuDAQbf4S98QeWxKb38S4w8gtJ+ZH+U+08kLrbmo9Jbg9
TuRyz2oaDXwVigZXZc7SHKQUWnNLZaYtgA+/ELBe6uxXm4/d5tkcEiX9yIIbRjSMHcXUTtudMDHz
YFgvrNKnr6ECwoFlprgROuXvh8vNW5cYQxRd5iql9Zp7nfz+6V1f2DFkLRH3wxkIUoNdaDYokJDH
RXbqKX4KTC3G+IXMa12fI67bT7UAiNRPnewY5wWaL6emk5BYekwfGq3PSXn7cMg7yLP4oZUIGn+V
kELjaB6JLqKQ7nw8LZkC2GqKGPeuOQYBkSOBaO0FA5iRSvBc2wpVLNp/igH4sH3cvM5F94Irx/TD
NNNJyQ5la6ZGR90V2SAGhgjVvmRbdBukrREEoqSm89OKXwThL9PJ06UB3oRRv6UaajBsctPDn5ne
ojMacZg7XoyCoj8lCyHRQmd6rD5i8Cak0MakSkj8nuOz58vG6pSzowKKFQrxhl9s8g0kwyzxbqZu
mVysUemnkBsfn3zRYYQPdw+zHmQpazVoFkEADPvVtlXvKam5w7ATzJ2TOOVvHxk6+qQu84BPjCf8
CkvbiIZpFJA4XjUeYJy2FCDoPHP6QsQ7+2WPqNTvqW1yPUC1UAy3RmhmUAlNe3zQyTYvITxymR3N
DMY7pN+8aed/WjYWdkRBqBDa1vUNL78CVhXjwSugY2qp/LviVezzOIOQBySupL9Ddkc6IQSt7+wY
XqkF2GZfnhQF9jv6dWdkOQlbX0N/b1Ik2w0psvCS22qxJv2IC8ctnKzg/vXOPy5Loy3XaRQY6Bs3
orGoRF8JFjipugnOcuDx/efXj6OYUoz9tj7NWeUZyEnqKjTp1ZhWiM4p5MpQeXznXZlDUtdDgBQG
yZ88eaDV76foMzBaQhirOHuMKERBW/vz2Z0Iq5Hb1Wc/9Wuoe8dDGs9ziR5zWc0senm4wrI63HaK
rmJRuG3uhjcu8EUKfv6hOabttlJJcM0EufDqyju/C69t6HEpe6hq0FdTCMHM/P43kEvUPWGcYGjh
4YR5onWXrceItd18uGGppjrAxsHz4no53FFOxtdC3FGazoFV9bfkqQlbLTuYGGUQKeslmxpQx0yY
yBqC/+D/RarU5bmKYwEXZOOs3Jk+ThvZv5Q4wFsT6Fzg35JspnRk8uY0B13GJoTStm79k4IcOfwU
aVokp0McUkIyFxKqCjYE7F5qHkuFRTLVdEXs0u0aUG5O9T26NiqRYHdkXfpLf75bBzhmg/J2dgNe
khKMBO2pc6RIdLp6CXmCOeZjmaPon8wLknXKWn/XzmfszAScvi94KLnU2PhZQbsz7V0F/eNaeIx0
1kxPTAwYzUz5wiaOPUKb0aBC3ZuoRfNICwmnvWMgTBdZb3dWNOpwhP01HyGhjg6q0CY28YGP3Mb0
HLcvlJ1FV/h7foQvQQSJNxluti1VbF1NWMEWSz2C23Inz8duBvIpU94nI78hS+fQv0b57QNSZ0Hb
srGbur/vokCbhNJE4O0apDCGmYXNWCs+NENc28BG8QzVSpT3+lyEDyM1grKKBkAhDaDoOUkoJnTl
N/heezc8pPMQFb5LUrym0b2JkQHV7ecycOT1JbV9865VYoPjZnL73FU2wuGfVesbPvbPMC/y2z2M
fHXu58nLmnLi8IDU9QnyNFmVre0BhrLflj7qCwldFO/gxkmAenlT2HZN5mKA6CFX2upSlILNmRh7
RvdMEIx6FOAs1wbgyrwHH/Kqsi23hI8JfRgyaZ2GDtjuXMREUm+qoBGQydcJgPfPbHvMNoYxQCyC
FixaED2mPgOhiuDBdCmkLckVpRrOF+m1vQWGyAJsf5U1OOEkOOfB5OxWvr7l/LeX6ZBGUDJMN8cr
i1HyYNRYiryTiyincn3GMKwyZGLz4ZuVgCZqkWiIZtp4pFWaHtDiwHf6p8wCx1i1TbrMdYwawntA
2bj9SMLhuvrrLh8dJkNZw2/6tDTHPEUMK7/3YqvMn4SR6GVeVThnbKxxh9cgTfleaz7ZQkN/t4zq
coBYRBCv18RexK7uWz7huMudhPyGYobaRnEAdXcXYSevwvLehgJObKc2WjvcrVzWUoDfhXVPVkWu
EIBG6zkz8BLnpbTd9Ua1IL42b4WogswzSvj0NWTXHxpaace+ld2gkapQD6eboYTNo7umUNE4A0LI
rkELWXmsbKMzmN4LothaDr0Rho8cWO0CNgfHO348Kd4/KJPnlVQxc5npaT+bmmfKiJVPt25puID6
aMqi/SPkTz7feYpcYn6UAQ+Su+/6TXhIMp1UKuK1L3wnQXUa4+apj6+kW56h6MCHG+RL5fSmZ7/o
LPsapapb++gQbaG+4cTf/aQAx5u6L2jS0aFQz/b4EHD1FHIi7oL/RiVCI3HInfO+w2+jMnCuRj0a
Bj4ESynmSkpeszpqJPo1YxaJZOzR/0Qfe6MULbBnfF3WFwo0oCWGLNgUIwVUpvtanjvX9GWpqmY5
8Re1TX9Lz712hUQMYBZxifPkC0pVbYqVN399BljGNGlZjdTZGwulXKMLCllRAJLH4OSOz1ienlV6
8uLd+G5uKtV+JJqDulJWPgKMxP+dxTddFhoU1/nVQS2N9q7c0fYp7Q0ZEYerEFtmseg0V7Tv6May
pbWe8EbLcClnRdGC+Lr2aFE5UmaxRijgKYLjiRqdns7WRi0bX6Mo/+CpVFrfpf/cPMcnNeFIeEvX
jTSCn6btJ7m/Cjq0PKoeFJtKzFIFsN3wVDXQuw8gYJ26egJfq0hBk18h+CsXF+BNZzqafsa7u7Qc
yHYRdfksOzQUHATbx3VRe2c/1rdRGi2E/wwv+38xO52f2QM9CCyAfgZrQn3ne9rwbQIatGy/tT9r
MMCXuaLfQhCo6D+Rx5U3TkPZ3kv6r63Wj5EQNrZvfh/ruxAYAcS820zso+EDmMQ+5+8Acaq6rVpB
XOG4mPmEpcQZW7rOT4O6unQ4FDLQC4mxln3X2l6NMF657VoxM0/aVsM4bT93lNB4bAr8PzUK8T+A
IyzksUNvU37OzHX2s5z9dNY1qVhKMkVPD77x232n0nhTB4YWzQJrqFcxUhvf2uIoZvF3D2rWpaHa
eGDTyhdFSSPqvHi/7olCHIvGF1qKbq514W9g2Q5Cw8AL803zSozgAf7RlCx7ydrCEk6o5Fh+3oL4
69hPvQgRt07gmU5CW7HC6NW4CcvvCySoJGCje3DKqZxuYoRjr/+FlS7ERwq0gzlxizzZwLtk3djX
y/UXuUOv/qOPMVCJjHjCr3U+67YGhwjJ6saSYwb23mtJVg6ZCcxYUImvodgvYfCnLbG3xpgqx3lG
J26CE9dQK7Vx6aDbJFLawg7nGiX/ZesXc0MGxh0mZ21hXcUd9aFmeMRIQOITsf0+MQ8sVxRcLsGl
XQLhxvkSMK/0T9KpqXhsc5EfAOulMUxTvVr209TkEHSFR9ue4cOUke63IFdRP7cOj2M88ZnXHk8b
NPuj11A2+XBG2Zm548iuG84XIS9NGNEAnDOx7QBmeCp4vJGCU7xpDffEfMDXrgEaASt1wd2xkjoG
0IuAhcFueQRIg8a4d+eqvUnu3Vc7uNhBvKtafLhmOXYXasmSotNsNwPU18dR2HI06nH3zTfe6f75
JJv2qVE7sK516HLuhIsZqN6/GU821MpLT8INPE9MZMffL1d/WwwDmVLa92HqDVp3VVKDODwJp6mc
6rqar8KiIpr/0noOOiU+gXKMuIUAY2h8AKbfYgTu8q3BReuTCKdoDA9xQROyKwE9fw/c0u9JjoGF
ZZUFH34aoh7ZU3OVOyzEpLKPqe1t4hHLDj6lLh3ErTekElTWtf40ndEOixSUGdP+KnM96SmSqOxt
KunqUNLngOFFO9D6/PvzW1feOSuv/H/Y2QzarUatqsUb36KYuPNlJcAppgCQZj97PfyDOJHkBqf4
2zyCFvgXjLRwO0vs8eM6b0F/no8mh3KKtt9+c/csdawPuVxspDNwvU/JvrH4eeAhoNbNOCZReGhi
fWEAvGLjHbptMPL3F+8OpIazLwYKYHJvnp4btr28BhF5lWrxMl1NIPivJbfE0IS19J7EzUC+LOVI
1xNar4th6KO4Pd+tMNu/LxtduCIXoreSOPZ9dt335ICUOzNPa726oVc+qieB2+1eAemwvHqIwxJD
yUwi0UWB6CLQ+BFMyUaYOxupMDhYGKKO58qDmSyRGY0RuKhkoq9nyjio9uZLd6FolmhG65pRodEb
KIXeHoElpPHDjAMEtMrDb5eVMGih01vGwTV1kPUhnUkxPon3YUXDAvLAPklR8R5vSKgugDs8QGtV
i5Z5rR66IJRP8pMSeL9Y9l+vX83mzeI/hNX8ZH3U13uVuA+D75TdyL3tGm1fTzSNlTNe+eO5VGdt
kEn8IhHCv/OcKYlSSCZbOYk4tYxCYSeJ9+vqIWV31+2dp49MeOTflyMOsfhivPrnVY+r46wIkaNg
6ad4DC/FKX8EGw6tGefarhOh4Vo90XiCP6qolWD5p3iUdbprQ4feOWTMdWIipGjEzmvWITW3Mewy
UAmZ7twERbd0g/ItwfQJF0ogR2bJzeqPw1TRS6EynwRVWfHBul3efubTqnfc+SqrER7qBwwBP0+J
k2d1/wOxqySe0ma8Fw8TJuc5K/TJYAT86OCJSWriNyU5VluzjQqCPFFO+NzJ5iBGdI4suXfKUd6m
zkpg1F+MmPe4vX3HOfNMPbfl/YKen15R1DVXTbl/86vW5UL2NljLEsXaPTyUEb0d/bvkP9oFWYFO
Qn4eaPiK/hkUOksq6SMMVsRW6iijf08PO40FlSJougJRxJTa6BFI6sDcWP8+17B5fmO9EDTPbFf5
5XgCR7VuUDXFTRdVpH5V5Kkmj9BY0WyudBtSj4oYJzFxgBgkbf1h3qPxkoJbmSE4nP2iw/8BMHR+
nAZChJXr5K61bjQDyChXo6lwgw0+lGfmwYM7TzRM5Eye+PpsHrFcWr1TmL17pkB8BhoMM0VSnZeJ
PGif5nUfOJUp4B8h1N0N3nGEleRNczEQi2LQTMm0yonmLY9NBG1bgv2RRiHiewf+wnBMinDYwY3v
oARP949OGG6ZpO6AdT5GtcamcrbDBO3CueG/K6g=
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CupVrRDHZjV2NAMUKyZqaf+H+qduH05WvWyKTnhg64sHsPS6zyae6UN8w5w7R80rZnJk/G3oBGIW
QavhosNCxWHfAKtNnagOLACOBoBtOC7W9NZQnLPQrebKX2Le1Z1jlWjURTkhfMLVVUvF43OV2AZr
jtEH7fXw8Qx4yfIdwyHCCgxuSj8+84rif0CrLObKPwjmced7fHljxtpU5khVFKxHDB7BiKLGEzQR
S6hYWDz/eJqmUveroNDRLtkgw+wChSKCoA63IlAFagcIdapbRIIwj/i6INH0OBwQd3J/IDJiCWzc
KuwSO3QlaLwA3k2+IDlVXIW5qmropb+FnY97UQ==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
HIJXVYD5wB3vfkwpd7YT4JZSzgRHseQsdfzPLInWtZHLB2oLpHerSWa+qbTePzeJuPXgKVwVUCcO
IV9J7jwYWA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
obl1tc/cnC3J4CpPh3E1uSeHIwXs8BBZI8SO8IiWVXwbWcsl9oodlrj5YHn+96D8d/7JROyfZlzV
h8LdrZq7bbnKBa1lYptYtRr6Hrk8xQabmCkdfm31DQJrSY4y/ELawZzZ0I9JHwtzrfEwlkGxIyFP
7wEW+oH4lqUGP+nJXm0=

`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DEzZTJHrX78KidN0uCM0AcRm0JC4mWk4fmVnMoYmnpifIfGGGqCn0rcYqAiPbYhbEozuP6nre5pK
bg7C7Np5s4tiiv9PamiFAVFeVn93AfAvcgUgzDmBDNsutW61XFx0hjacg31PrfUx5i/pNrMfenNu
a2+yGIs93adl3+Uh+/M=

`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LwxxdZTZIgUp3Kzbxt48kG/96WKDY17q4wiCvS4FqLsf9CB+fUSkdAuv01U5QFbluzv/kOMm6jZd
E9i98GRFHCwWvqnZHFa6/7lnO9f+AImPv3MJ781NafroifGLaeUb0yotRG/bnbIh8lOQODry2Nlz
M3oicuoLw3iof9JZMPLKT3+Zqx+fN2B0OFKD/5sVOomcfJSKbZaRj9i5s2Ht+rWU3Q9Rp6W4pzb+
c06Juqqqc8N6qrCcS0Cq2g6Ty9PGDAxd1apExzCwLCDWSJjcm2Obrz1SbBLBdNbkDa3xfZzwdaPw
rs0YtSnWSuHzDQQCWrd3VKZrNCws5WsY+h0pNw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 148320)
`pragma protect data_block
26CAXv+bB6Jheg40iBuGQerL3wR50a5yhYO7vCU/edluH8l/BVByeJM+MUmTudTYMUgdDYBZzUdP
DWPvV9wkNHK2bMlYZMAVRhCIjpIuvzs5GjBi1w869tComAvMrWCV6aGiIDKLn5Eop7hXriUjbCbE
W5C/5ChjRUT0Br0ucfxJjI/sRJj4bjrir0FqAGP3/FA2NTnIf1lTcOg4b3OdSmw+hjvmPlXFKSYJ
/9LeSQoKgKJqh8pgmhB5swNKbnKu9vbXSYUE8dEo6GWiKEmmI2EZqCph/axIhdvclG84rXrbpQnG
JPpDPjC5cy98Ww4fXxklXZvA7JsnFb2QdEYtDGVBGt8Ks3BzKmz7FcqlQqycs9jOZ+lCG/zbHTDi
fvxApL3+D5kioXiQ7gbCITIyiVZePwfUYmr+UawOsenHvtroJWopaWucCKAowQOtCVmp7DpTBDIK
NC9coXGVi+gZkJ4XholDtjaYKcIaClplJGZNzMBSc7CBJnjm9IAXB+4jfNLDyjSQYIb8lxCrVCTy
HlGbkJeocrvjOcFSpxvWmQMQscMrtVHpB4jnmiDaIwKA97oQx9xTea1PlbR9UoDHao/6vsB8xFxw
/2JJMPql9IztlrLOdL2q3pX97NVVUE3jbFkWcq3f69yFD2hvtQt+MmrnW5zq436IXV+uFcc65A6H
lfKnVAydOEBjDxzJ1buF/cUl3Q+byn6yAJo+S6Is2wmt1kc4oqzFE76rg17o0IKf/szvfvBw/ClL
FZtp+uaoX8ZOgC9TT900sBX2GkVT7VzwlVOMAX0LnTnkY1ArwSHOpokXGeDKBJzSHPLDn4DzEY3+
sc0wi+5dzeQbFCtdvZjhkZQzFXQ/0HxjqAHDfO7Rtv4j4/imvoR1V2cCAShQ89daWwMZ6aM3UdJw
UShLab3ze/DPCWqcRCvzuj6QCXvGstTgBJi4OrEPe2kBu60xm/xl0xv357O7JgfGq4wavsW3Pdjt
Nl8XZeH/BiYNhmKaMVFfdMX/niqiRrjgxzyNPEDsUu2OZ+5er/ajxk86Z21sYs2JuaoWLILb9IU5
ppxfTYyuMI8IhI3m+4p/V4zRn6Q82ITpVWATfynC/Ria3upQfe+wBu/fpJkUW8C5Gz2/bx9VE2m1
ay2O8OA2HXH+SoX3+ok0oMpNmlL5ptG6MDry7KWXOGtYbb0S/P3K+gelrsypjFSL5vtpUQiwoGqf
1NO0TYoG9hJsQNFmdF+CLKLZcPrxA0IiwYNGk4pFRSueNryh95+RkgKT4MrcFgGm8vbsimHxxi6P
dtWfBhzuj1FXtfq7NA7HvOs2PeXzIlhosym2Mcst4ru1nERuFIx1YQZcTPQxhUnlUZcoJqNbDEhE
yzec2OF0TdCswdyWaItNH0zscQPX0T/QSBYeS5fXQbkshH+NV1NhagKbiPR+e6NdBwlCUzlSz8FQ
NyKrOu75jl5smIpl71kSrZ1SDb6x0be9YuTdoliM3SnSm2h3ybYIr+ymg56ksk0hTgYD1dlmKlLr
2Mx/2LHvTTm4JwznNnoN1c4mJn8GksTz6Sk8kqGKgKTUHiwxQ3vv2Vjs1DBWDxa91oPilTgkK8lr
6J1zxOPHPJs9fmm+FgUKzuODVVVqQChz6naCIfuTzB5xyNXBnd+O6dRmwv/Kd5QmlO0lp7eK9cEm
7YzU1SCY3V52HQb7WVreOjSM2O41W0ybBLBUAgolrbigzYYwQzguolJ1Btoh7weoRXlJwuIWpciD
Wcf1zfoIQ1Ih198BvFru+GkKzf4ezjVS39DXdv9sSPkpQ9EW8U/O3HAGtuhjhgJosGIsZULaisQs
4fygGIb9vU8jFHGnAizizbhgjd6/qZHD+PRRzgcgq9gGLQC+Gss2ZLDmrofKN7xN4Sh/DflDW1GK
dkv+ITln5llhKaIGZcqcm+LDVT3UBZbE0mGG29LHXFHxrPRNvkANn6Pltcd3egckTy7R6kvKpK3N
Vd/oMPKRA9FwZo+Aa1tFAM5SwadMG4ZOKHsZz9CCBz3Ai3MLXDUJ7go7vtULZ4xqjeJgdEMSe/NM
Yf1FOrhh2ZHiBECZTbx4Vo7jAtDpR573ra3HPcFiz6+B1tWQKmGiOBAlW/sJ0K4TY2IQAECksgsQ
OD5zwHENV62xZBKeGyTGOgr0CenCJHhVy1rO4bqU5F9VlrpfcOGUKyiaM4FUUPA2W9A/fsfZJ8s8
MaCBgDDKzezN/VimVI6EQ2E05nOrzbucOsQTA/KOiRN380znQNarwS8t3kQIZUadu/9WyjPuMcI5
dCHRv9i3FNe1Ik0dE9t7sAXa7Ktz314bMraI0qbn+Bm/UnSeOdw8ESYqAi+dgRGL/aOUsf4V5Ny7
2OT2+PNZyu3wJQrYHYTv7ljoJlHAYfoRr/fruxMsq2g6f3NRkSUEusu0GySVg5HEG2gnjq0yl6Mc
IF8Mgjh0qB9N1aelemzMlab853qcC65Tfr0lYhLMR7e8L7rH1J7IF2MaIqc7O9hbvH+kHluxevAe
ruahHWygq4VlsG0obba0w1KtEFWm+HXSwaZ69PDpNI+oQegJgUWH+mN0EpOK6CP0Gsjcm2G9N+Zi
+Rqz+sx3lyhg8gjSZ49X5zCdR2b0CJgOGNxAfDV905mC5+bqX+TU26oIJ4pWoqbzm0FMX5Asq+AI
/M1VuQsB6gnHchlWiAg8qK66w2mZKMea7W/eh9SARta0VrRYCod6MV/umOazTTixm70B0yvzOnL2
A44Og/NSknCmERQmFN0/uIV2m/fTlTBMzlZFJ7FYrB03WQ+izYdI9RJKJSPDJNk0RVHLwr8kSLPL
xlJUKkEOhZVLnVHMn2FPwwZ3kLp9FNq2yWEA1YZCoS07ysjTwTMDitmNgE4UvgJVXxgLsiN9fWQF
csg6gyKGfdAy3RgkbsdRnvi3BO6pE0UhDdyHwcUcDrx0m1UcsLwxzyet47jpJi25rzzmNF9vRdKl
XyILA20GOBJhJA6QLGuqm/u1sJ7BnqKNoBNLq+Klt6FQv04T1Jz5IZlC3fmQsyzCBfcIyPr1wVPt
CiVjFAlu83F3QJX6i4YNbPl28wOqaWM1wFTRpc4523iT0nO+mzfHp7iXpV8yhfktwspRqUy/e51/
VVXFX7aZ7rMHaEMMeIPV/ZuaQblcxbwZvv9EZqxfxnLyMKdh6kQWrKednHaDsttpTQCpLX7pXrqb
llJqrLYICHLv12jupr79RNUDsjioHXMnpuHcEvkHS4lv6JL61E7TiqQvdYelHwV1Vkzen5XraNmK
ZBWmEif70JxxsQdjnuz/+mYpWIMQpqppZuPfcQtv+D1XjB+ipH7AuWBoInFC+gne2BDJhYacw4wZ
DtxwMABdbREsf3omnALAsAw3zfjDDLsFlL+aDJzGTK05OSMqesMjN/3OZXvQp6KZPFI7VhbAxJ1Y
qbOCv5futPE59zSS5aV8j+doLwtBmWYp/PbUF97PA+MLE3kA34/FwxPKdiGTLkNXzx8jBejmiv0E
lXg7VJpCMJorf6Gx5V83pCH904osffJy+sdn2PdMI3JnPXIgfUwmQ/MwNCRcslViZRZ9t97KZVM0
Ca0vlLYbAVCCAXoBjVuoq1g9fko56zpLLo+USHcwSmwXgNkKS+4MKOCyUbuwb7gxWMAKhnHpdvBH
n1Kf++/NAsck8ldnTCmgsXit2LjfhTmeodXYar0TciZJ0MMfHS3t1YJbiiBtRMNESMlOqMmxGuWn
3gb841586O8qfDKgX3kXCMSx22F1f3P6vYlaN8wj1GemVCU0kPWxAcGVJU7p9yugvw2y4APz+q5y
jxoMBwh/xYves4l/PEkUQXS21WxCu3+Kus/JKDdY03XFobigxFuA4pnWjT7ldAe8nzHTU3j/kwrA
q9avHwvGwcHvlOvHMUFaEEfcoZWxfVLJHKDXzXOCT3SLi0aSWSOugN79FGAe/sjkj1Wulqt03Vd5
12aRhSkWzbVY2aDfaXcVUbJRAy+r9f96gvlvC1FurlfgMV6RkMhPkjgNbzJEnCmrAb6uPN94SWSA
SMDWuxOyHL0BrLXv3xQ4Md0tS331+54Tga5OLwA/K9KBlxKY64oVF5ujYMCY2q7vUQnmOFgPxTCz
O0b4FyR+nQF+n/hF3om7yp5EWiQFuXTb05EBpNKD70gtqIwSlVJiG72unEEdvk1wrJcJqiAymN/n
XRU1b+8I5+/G4LHy/1+RjBdRJreA8hi/5arfU9EPUKT25jTuvEjROoQG71uAfMD5uZR8/S8uOxLL
q41/QktwodVrFAy9lM+VlZ6NqcYg+kQiRctFas13kvwu9q1thwblR4V0eYdM3jS3Vu4ueh9D9u4N
FhF0ful5EMAgI4uVuX+uCn8FGz8SFjwqIUtqNSJdBPsnXd0JQXwibzJ3B0MnFYEsqnxzltX/yVzu
XZdT1+aPGk2+hzMK/AKkBPaiEUUynPI/oeCXpoavvFCKARkuYGrZj4hcSPxO7YK9ZPZu+GfwT79G
+gltJhKapT1GObfsPNvYL/WyMlOI0XAR+JJ6Ns0lTUeyAiw1mBujwC9vAPkl8ZYk1941RR9MiqrK
cphOCAG26TPntMrNxrUsfGGESoAW+Dh+D5HftIhRSIJTCViKpZJmLw5rmOT/HTsFQNfc//SpaeJy
9ovnXUrOyjTOrd2aT1PyRNUwKBp215CQiL9IbPspa7KN2OXroRJoDUPV7G4W9jiLSJUXepXRS91C
YppiLcwaPI5vKb2Zm0VTmefDgMXXxm//E53wtl+koNbMGEEyqNIk7kiwvO1LmZg+warHB9ujHwnN
HRXGuc28zsry+x5nmCSEO3oXPd65/xW10MyZcPbZQOdiuWrhFxmcVQGRoi6oFmC3DqjfgDcdgpjv
+yZ7BB8A6j7Gj40Af+poGkD+qSUTgJWxVDdmaQb/L7UJsvMtvgXybIQpnhH4+HlKZ+K/Y7RfgvC7
ekH5fVTyO4QBDF8VQ2oV4RGHhexz2VBevEPP5ytFcCAOyBL5LTuWSQB5ocy/aSNn5mkeSe6Y2wdX
LsDs9DqQ6Lj3FTTjkVZZfRX6yg8wiTGZdFsZCoD/WrOEPSCropviNP6u/nB8uanAKnWdT/I+fNTy
6NyR4UroY4flyI6YGtXuPRi9tTMd4SYcSIPn7goGRX60cMQcgKrRwH68Ym76TQ5EWHMPGpGiCTDg
yxlj5tWKKVM8g9RiPVJlOhANSjjBbvvy65vtCB5FTtmkOPn9m2waVmOnU/kpvbW8rFfUyE9iV1cB
LByN9cHUzqkM2ev6wo1AullfdOQg5snKh4nhzjL83FYw/uDWaD12nqmqGqU8RI58xftB8G45WrJh
WnmGOuEsVEKsl4wbIXTEL+mOLHm33DVhtuzpBQW/YxsGHa5seUAQDyzpoI5R7GN6IG/ZP9oPAsPP
48DV+18o/OfLQ3DKy87SSElRR7gRH1RBLsJ17MT7IGPw+irleTr71C7LnPzpN4rGqb9zBe0oJzoq
l7/NLv+W17lorL7fNyJ1NJdUz3K4jGB8O0pJyzpXV7qizsWCwpB+Nb1jEhmAAqWw2L6s0n0CwJkz
93iJf6REND29CVmTwKL64XGt21o5wGyKiVFrYe4CZZ0hdA3/zKnxfQC93N60UT/fWWx/4u74yh2Z
oQxKzvkK+j6qjet0h8G3XWp+g4BYKVI7KpX1GCJ7edxTapzfclxBR/XuQkFbc9t5ZJdtwG+GFI8i
RihQxZRW30I9+4OxnTqG54xicZlldvfz7KNJKPuTojxEvEdAFVGIJwxvf135DG96PKLPE7M1jfaj
4I2exZR1Sr8uDFQ2XujwYsqV8wSaogFskgxJtQFY5HAUYaPdnzigwco25zUmyfEHmOOQdcy567p8
G30Vc0ClGPVxVj/kICBJ1ieIhDtOyeM+Ah4VGO8cbROU3dwdenhYjEtAAkQAndEPTupCS6ployN/
+qUpmIr2Oxg+Dv04+dng1kttBNonoE0mUQuRtx7QNtVV5Y5T6TsSJAbfta/QPARCniYcuR38EdDQ
vEXI/Tvjj1xxIx/0xGkGkLrJ9OiE5OBw26i93QiDUBS9cqTsP7vfozg1UvtMPrH+e41TXxnJRFFW
Xg8wYl0lvD/TVBdAdJVI37e7Vm3EoieNADJcxDhDIPsBRUhgXFYMHQvcu0Sl6hFsgAldkj4RgFmI
n7Ph8SlQ6JF2Xm0DSH+c9nYG46L7tdvl2c+1l3CDAtv2Ghmi7VmkfwgHdJUDowUAHG8iK40NuQi5
/h1WcQEiW1PgrzplEAfjyJ+lysJxE6Z8Uehkr/WuwAryu31alfchegDlg2a3MHGKHkwwBh6Xfb+V
h99runhTOb4chaHFw6flgMxA6veGKcFTOnCb7cfI06hlMMYhH3BQAWtYFBD6EPeCV+srQXk1p3Fy
v4aS8nSV6PQhS4+4/M7Zfvw9HgLy+k1sGKwx6snaEJfxo/waJR4b42MEZIeVJxZm2HpxEDKj3lFJ
kj/iZtZxVu2sp+E0QuL8f39qHf+EkOfi/eQLSRNGKA980n+yU4edHk5z4dXtU61eQ61zmjeEsXHa
O6LHzkqlNXJMogEpP0DMDCgGbtY5THKceEqic7T2FbTV3aCkkvy1X6tEhk4LP/vOOMIeQsYCg3gR
+ASWXg8rKAK0Pgk/XXt61B77Uy/puo3hKxwtApaELu+7moHcppX9MxXV2L0qvdbG4Fi0XO68V8dA
nV+EXa6tbbylzBM9oyzvTbLdV004qfOScJaOh6axvjOsRZouYmNe27l/Aq+VqXXN1qD/yQ52WMya
SO6cHcmIShpeueoidbCyZwRWR9+wwkM6dCI+kzkB7635hpH46tXimUdWzOYM74kBNVOXGQPw56ZW
b7DY+/SzgS6lap2UENVmaDkq0IG5njLME4aBxa8nnScWV7px4IUum5eXAByjkX+Htx9x7yIGsLry
U/Cvcr/AkmLxqp6x9YoOTdO2On1H6yjSbv7JFho6NfUhjVI3WcFtf4OPqY9Rb4qu3VmfSOwXWkAu
nF3NpmRQ40O6MqPt+/UFsey1t9aaFO2/JGTKloEt2yG63TdSTpABnGARI6/6HUmn4Ted1BdCW5/F
pd6MDP/ChlJ+w/R9beMOy3/oWfc+Vh6nOueG/0p0c5otDTsp+FieJGfHg6m59c6sJy/An2433ys8
u7FF+bXs21JMlqDeU9Oh6N1e/lUfIk/yE78qwJSwxwNHCiwQYnbm+8zxv1b53nwtve1e2pRgaMmX
BctFW8ktWFFFqVkVaNWYVEevqdH7koHPpSFCosAPdQtF/gNZ9866/iU8GdsDemnQ53XOXBfjZql0
8frDmnAUI1gO34YBC/CTmt85juA1VgpABJu/H1tOEa6iKqcGGLZ1/8Ow7b1wAMYmZclSs/X25wKS
uvzrLfnNPceGh5pbMDOWkDUp0Sj0pyi1PvaMys14HxvVFpx8zboTjwHU5cs7sojPN/IuVZT0L8gs
3Nqvr+Il7Il5OZYOggePtugAZX41MYCQ2qgPcEHCue7W2gccCjHV5DnuLC7C6/qpuC9o26vKtlN4
ljON0bWxA50fcCL236WW0Fghi15ZOBqQjzmTuoB4g+s2+kQlQwtE0WN5eANFkGTQdFxJ8wit/lo2
Qp5yUHfHs4WdWsVv/cWWV2RGYG/mdpiulhJ7qNGqofZ+lZ552Oy+h6mvNWiNMDaaEkXqxJVTeSQW
aZbBcRumrbTbVORxfIee3NEQgbW6R9jChBQQ/EGBRMyhZHjECNuO9o7PgAPMZf9SSTM9GRlVP/tv
Afi2/EzNGHMXV/J14k+g9Zf9NSZ4mNdStabFdYVtZkNfn2OtTj9TOZDxCxtdFuZ/5HmnfkeQBKHE
CRGymnIGhjuaqPulRNGA8PwmMRN7fe2RwqYlmiJx54nk9gcRSb8WR4WRevmh7Sfiv2oHuHrE7mPP
V7XVQ0PlacMXwtMAgvjYn0rQaRaf7a43GeaPbimR3YwDv1BzlDVbOgo7OkG1O5x0CZ4mk+x7dTaa
4Ace+uPphxJ5OhZhmyZ4XQnfp4NkKDfvycci/zGh6Rzeopct7xbXdDTBZ8YNiNouC6Oe9EsiUCQ5
L4QT1eQxZjOCqKcRlqv9InZn0r91YHWmTfS3RKUSt4iHKDVPhPrnvSA3B/mtxgdTwpE9Mucd1h3x
iuYbLph0AOw8iuGV58OM92mWMrtfY1g1h/6Be3qEtSReYdLIdb5b3OWs4/HSvXSC5zbTDVeJt6f8
x1gZGKcw7FH4685qXj5y2hfRgM3kOi8WE4XMx11T/bkpZ4xNqBZfhRsWWI1fPXz93gAqGkaJ2LQH
YQg47keSY3ORWpky7YUwLCEOmEiZHvJ8L0+UmEs3OnTxpulYDF57ohKXMRgXQENYo88DUqX+YPSM
+jNSVyXM9Awhu50iNL98c2HkbJu2M7lCmUqzbM92HNbvMOfxa57YPgRsXzjIWqVY/JKHpZLKw7PL
ifK/jWV1+UGEHP8f3qhB8Gxr2nluCMUTcjrt2f8HpYy8+VZNpUwKn2n+pJ+HfXtyQPv8p0nJaEtG
Y0D75Qbm2uPXz1ZBIOpqso5PVJqJ1zLj1OgsJFZjc7j0VJIJbokM4l+Ybi9RU3J/ZRHzFWI+UsZ9
EGdmo8r79puvVoFHRB+3IK/P2ndZlUENugyD0MjLOVO95yD0FTUHfkjjzS8RbAFpVRNVjxM4bEfM
ZBufphy2mMu7g76cqttmTROcwps9Qd5Z8V8SBssD52P6SAhezdJBtidfK6/dtpm6cddPMV/0E5nR
dqMNxcJB4ffCksMDMZspIvBZmWY/XYvJBwwpDEGovrgjgMERD4ac5/lisrunpEj72/nYuOoGMVeK
ODoabVugojcqP8aSvatWTsS/QN3PcMgV1iW20y/V0wELrAhTQWwxfZpbFQacCDalwuSyTW7QPeNI
P2gDQL9AYnesLUnCoso5KJs27OUs/vRoxQyCMu2yowHRt2B4Ig3JAZ88XgM3M+InQ1JcIY/EpQFr
kLjlF0ZOLeyZcaL2d23+pPxj/zmqu0Bl9VQ85ivaDTzKEiZn0yFFABFLyF0TrU/cZs5O2uWFWm9p
UgwqAU5pKe2Edq+rmHMvoJuS4i1MI2aDkNrr714fIG0dVeq+elZ7JS6B0+nAnUMsGabtWC2l55xE
c1EY/HoVgjQGEK2oYMf+dI7GtXoC4GedFC2SkDv0HWZv3ft9Sr6OW2ogkgKR6l5lIblGpi4fTBNt
PcFglb3V06JilH7faf419w2Ay5S3kJSoh+wJofmdzF5b54Ji1H9M0wRQZcJmnl/5dm0ioK9vcatP
Ui/AlYhsuXObbM5PQ3PhvCijj50Q6ThtUK5/FhV7kqk08L3G9Ujr+XpVxHeXBY0XTNBYDKm7mx8i
RJdhkALNbxAGcQy2TTA+WzsSEaY+TmEkhy078BnRDHTeGhqgi0LvMOS7tpQIN87uzPcJMV0PvFZU
L6pwnvySnNzonQPy2431zhHfIzJGa4np4Ea2mjfxHKJDno8mwwIUqv0mgUZXkZnu7wXkaHPY/BwX
cV321BXAQAW8MbRwWeCZ+hCpDQ++Dmrz5x3mdzHJGP5FEGoEIDVDOcUg3e42aokA79dMe0rVXOeY
QtovPETfLzvQfQwBP2Q7U7H9whj3jYrgtm7MJ3yqoxh2lo7w/bR48X8xPPaTILiBMucAeA1NJlR5
HEMPMczef+h3b14A3ijwqIDMbJR0fJLiTTJWUHo2tA69SKZotUWjT2+j0Tv+My8dQNcdxUWPTLo6
o7PN5XXyJKe9xw+mWecei5kfIlsJj/fDg+rpaLi01v020WkiAffAqZ0TsikiLBnNzF9VKpCP2qvz
6Sc8vzpJjZlaIk52IW9xaMMC+PVAAWXPs7oKdLoSlGkXZCLVHGq0PipsC00e+Vbc4AGLMICQMyZX
eTIQErjCBrEG9fJWu3HxpBx+gYe00QSYxSvcb3dDrlOlBlHGhnIYTl94YseQ30vpnRxLsL5nnmA9
wfc5ZdkZLz4eVmxXZATqGF1UA1nVx56HpKtOBDLcnvpmQqOmbt5AK/nbPR5JqDlZf3jiKl1SOD+x
zYDR+g/C8FCN/EExr5Aby4mmE7maCQNMd0CXmXQiKShAQG3Hpa3XCfyORVzTXmlLg+hKVVJVtxOG
LocJTmPuXOETgzEv5BZagOGz14Tzcr9/icQhnALl0xLRwO0xoIFfePhHEVLkjq5qFP81WA8lwKIP
OCstXTF0XYQ//qUfh5HuBi5/ZoGIUwDKz96R6Nbo7fwsMRAGXSO9V3L1Bs1ZsTSatE2f7NNe5gMR
H1dRaypCS3MbzbaZxzZoDIxAPM9dAKc9RuvKGUgiKAkDi27JxDyEcCd4zS7VaWSxQ570zn17WMbD
DnqF6FwjaKvv0EDcqYETlbK4tiFvZw6r98DMHpRR9bp78xmP/pwD5Z+OYsxffVEN7+KySau7k0t+
M9omYN/ijEGT3lMp8IH2O0D5qoQXFHgLgJBCXjRit01ikae0Lj8KYkN2eXgPoVz2kT6LE92en8dV
vw4PWumsLvAoPhVmxcQNfYEkNaCUZZDzvYLUY7pScO1g62jCh8RsXW026U2QR5wMqr4CbdC3OlHm
B71QlxyZN3p4bYHMcUvBuMP9Tqr5Xd+kmdor1L/jascSmTy+CLC8+yf5vYRUvdtdvImqRfpfoJVe
HCHwQkUgeiiFxmAkX4WGHT6QQQjGZbn2cj8WinHb43Nfiuf9WMPYD09T9mqoZRv2+HmfonWg2RBv
OIrqVm6kFa4tmzqRSW6haV9ienN4O1dDlwuy7rruUznLdTSAh7q7Kw9pPZzZGc12JOCLVW4uqxTQ
gKKDQ95zzrwe3jLdmbTVipqF6Ibt2mGKWUXkRsDkCSw3HRPELEIK+Hn7ienv0lBsDdYaau5PgGMA
su+czzNwhtN4cyKppvRR+eUJ2izEaD3F5KwgNTDcUPZfyLrZ3w+u0Le/QVaumrIazM4YiK+EyJuR
Sq8wwaIDTKJXc+ODZiO6QXhoRkZYm3E+0Iib+3NkSS9CJ4GzfrE7dtP61jrYUAIOGg5puf15fvDN
B6hWaSBvhKna/jIxP7PtrxqTpiLKgNtEG5np/kw6Xmcm+gHmfHCH7csVu0AOYvGDN7i0LXcZaCmJ
I4OkzBNBu7TOtpkqZrHtOjY9k1aWNmT2iHEgaNFfrsYXXo4LIGUgMKzv5UgRCERNcf861LQ3YfZL
ycDBmo4PKuIwnkzcVhYg54Cr1x6m6GYaC4+p+hA9hBZ0xNbvEYyxu7DWsGia6T4h5GRyd7MvFpdG
IuKAXAdpedAUcjOUyiRVL1OneU82nbLwP4Yw3sM4s8s02hR/lhrDtT7u8t87ad22O1/6KV41ul48
jP36P8Etkw9FMX5ZP1RWsm9xsmdtP74TCgdTx9OdomYF61QrW8g+X+QVQImPtBEClN60G6makgge
Y83p3+WgvFLRZk698BSRM2WO087Q/N43OPbXIKBQw2TYgUk0PihBjheF6dq+R5zuoSJxzSQL+hAt
85vejImKezkbmEAAxDNGEtU89bp3NYiY9ffNyZKz3RVrPhHI2p6XdNY8ftvyn+1E7J10gAKZTWHT
7G4EO48BYIiVOH7Wa8PDR5r2WfPjyQpsEyJxb5wIlrPKy6fKaKQUP04EFL+Ia+n8Z+T5hhiw8vAc
bmyKs6fn7abkANt3t5AqfpIMYmI6vzV8GYJrV1U+ydNen+p5hTpJS8wpOb9E6ltmoivXsT8inOvQ
UdciTOltV9Xz3eR12b19jf+zX61SisGqMjjIjPQxwmT3oatfVouE+XxKzwFQkmXuDWoBnmKTzgm9
gwOO4GGVmI4Q0H1WLmv3Bk10l+rL7WSHrHcvVjXcIH9FlPEpShzReA0i8C8cXk5M3Hm46TRwzJ4t
CRYvTiEU/NZAdQ0+rfp1An3H/sBMngGxg77k1JCCjHRLg8kGY1pUI2BMhVl9MSN7cKZUWLptsatw
mnnRCyyH5EYAGisKt1AuLCTYAp/D0pJZ5QyhaubIz0TDkkVzXfCajyyjiJoJgVwC5CFxOwjQSk0E
OsUpqy6fulobOqwlZAXp+MOsUj8GIKhz8greFg3zlZzcDM23El9mjrGkqbFTgoUUX5RETxI1C1Ok
VxmHI0rPapMWC0jbkuOZdpJ3SjiayJsfWZ4srgAmx+uv3uuacpo+IZwyEVzOOqy6i5CI3Tpe6s/s
tN/GK6JvugPvRUSwkKRjoE8RagJohPKmFAZU1NRkk5Zzw2RVnGzKyywGvD6xzVRWMalPHue5zwFl
B4NgLRhTcjjh4wWrISwixA4vm+Flq6MEStr5qcc/9Q8Jnx/EpwpxllsE5tz4OM8ta/jgQQKmrDHa
4wjPavRvOUCJAQQVmJPi+A0lHVxuGxIOoHLYTB/l3VWh142fPqKob9PK6OawJ46Tj7LwMAtyq4Ou
zJ+h2hpG/0Lzazg5ouN9h3ymg2q1Sxj0fFSyfS9qOEldHXJcMnf0va76lsFuTK9e+KXcroDrYJ5u
cI5UFAh/jQpfFpOv2k86zukzLLUKR3/h5XNO5P5/bv8Fhvi9l5lNYl7aBE5l6nVsCGju7ZO4XuQf
LeztIBmnCek3bhoDI+jw/PYd85rcCGe0vDpQB0aKoM8lLgN8FFdoDslnqEVqdtxxcbgw81Hd+8Si
nYRHIxAyVb4YJnhJWpDUDPzNkkHVYS5W21T0+e8NvDQ7ykoJBVkf0YRqvq1Aupru3GuQCif2cOCQ
B78xl4TmVEV+IyM5a/6WAzhtRuJp6I8UwRK6xi9fRGNb7Rli6n0B/O6xI0M0OEuXn5Y4VQOpz5cr
k7AYR/hRvtBRoAT1ZGaRwRoHiEAggGN86kczqBokkos8ZvYAWxiRZErKuyUC6Lm756DACUyRLwb/
dQsPDWz+XOoYsP6lPPCdwuHffjvrAYcy8oeKLFnjQWqb2elJU5ahRjEoXlSHjyxTxqm0uTSTSscu
IPZqm+bVEOhAittTsSX+emVKxGW0unMmmQNQpOyMj1WZ7ljx2IDO2U/tpA0BJkReAWeGU1+bBu0C
wBnhJeqII+MrSNMbTq72wLIOo8XFT1PSH25XXyKagDQ8BFlZ4txCPdcPaftbTDxG12LyOx6JmedL
XLP6T3YU34ltwVAbsVlnrrrNf/xE4tEQiQV9ZKgL6rqKdIruSaJvb/uX3OV/lg5+VtI4phj6/YPK
b0Rtx8eObQkYapDEhEMG3vw1saWqPNCY0nOwnnQs65pVBMFE0hGmDzN26PAjcl7qvoWVisXVtQE7
TU/oeK98VfeFWNo3WKLbThwYT9XAjneCz53NTvqnXbunC69rhlJfXHDNHvRaJ3cUI9YdL6laeOGM
jYBitggp/ijQrBaPq+6z3hxUGWeNxhrUePxjidQ7uyepwyeCKYQG1tlTbERQYImKCQr9MiXJhyzv
7sYfzB/U5IxiGWlXFKTB+Un77LKXF5vHjf47n5h0Nzc8CvC58P3NPsWCf+EBT8SS1BMnAf4vgHaD
srubAJ0LZSvYfP7DcNtm54Qb6mzIrfVjdFR0fdRkE/cidkBuhwa7iwUPq4BdkN2xD6+l3pkCnAx5
yWxa+gXnHQmYw+iivfuTS3/ArnjMBvfc9vzyWtm0cH8nOXq2ij4BTOhf/cpIQX3sYv1gJXGEgiJo
v5ycwVNQqdIkpLGtavbCOo9Ao4CrKYvQ7ePOfdAcE0a9h/yiNaNSaZ+aFMrAoqHlWl9h5i5oSIWo
gxUJxoCDi6TyyxCsn8thVhiY65dPM6mi7Z5ByPTtI/0jJLvLVY3KQVGa6LKqNHmxBQdSBzE6NL7D
ryEDZztJNRBkrqok/xM02ZyzG3DcRUp89QEdGO0slC2KmDtTox7scGhNBj2JqO+HY7nTVEJXD3FC
IKy8XKxRR/F8nGgnwZZn+KYnk36v+ccK4ng7QagYeCQfAclxjSr0qwE/fB6zFoYaDz2oBa2d0s3N
kqkMYwUSdUOTJGK6gPmJoBKSEeuPsqhqfPIh9YGZz4LLlQ0n838B8Nq/mJwmDMcThNu3iIVaLR2u
R+ZIzO1uqoLvfz5qV2a8PeuSUs66t254RZe7dH7U2c1+Xwga4Cl9qg78v3OqEP/Ilgz9W5ptQ0un
XbVznLnWkYvMAn/PyIIe5WhBGWMJbVcCSKZp6vmFx/LHBbX7Cg8jezrg1Rw+FXw3BNuYdO5I4izf
SG0UM8q5sxmBm5gYCUYlVmyk7OmSHmtrX6X3zWpSahFhCK/T8LAePJOyBAe8V4okGR49MxALQ1t7
kWKqi3XRI0t22YpYhOQyHB49k+IK2oBnoq/8y0Ge94F19/tk5ZlbqAr6ndDvzydeJOC3b5aGctvL
GteyTobPqo0WLaS6HlKNDAY4CoH39lhgtBcyGI74FXDvZNRaY/gvbzs9IaCICeRkfX4YGXdg4kyV
VIkGiStX9RNZ6SEtF9Q45bQxaIXo5KtWh6VgK1VhgVLVDcgnAC+VU6a5WSO3LZwyJngndPXY32Sv
7Q35xsmloQ1GRMReru2pbcv4BLcA1x0HdpV1CRUoSO33qG+ifj3K3uu9sMQL9FwmcPdTGpZJFfD2
jfoA4FCzxi9h3LcMZEZ3ifmIn8b92jihp/KJa5tAsZH+5xbvn73ut7Tpr9f7SM8RAd0zE1ftB8n8
99Mz1oi2qQAldyyH/C6WweS7a3MRkO4Yjm1erYW7w3W3Gy7Vhjp0u5CRXKcvaEh/uDutBZ56TZad
G0DFCmkx+9yxamThvkQ40vywBdbyv3oHiUBuqNsiQicGU0iqhoR54adcxNyEHvf34VfYTEgGMwij
k+e7ayRM+rdNsZKDiptZAJ6WiP5HnQXWsCr+RkDlG1jj4rhfN8Nl+DDlS93TQ1Hg4MAfXpcbg2Bi
BoSDHuBGN91Xl2bX4zJYJnkqMcIKJKwP5GLj/8opPaJlnHIBqdUDL26/JxWENDyjoKUjm1vI9V9Q
5+5zMG5MkxYTb7kGfsgoYrXLPJidDJuueNx/wsCTFc0L4QP+/zW1oAiG/nv+u6N3etudzneSt1yF
FEzQut+Nwtug6J238kWfs/HVNQny5QtZnNsPnoSEWQe/59TD8NAkdaymleoC9Hm5FJGjLWV/T6fB
0RMn3sVTJahHT3RYnECF0u6C3vMTmMgaD+Ah0teNIqKxknOgQ1IYtyCEqu7VSH8dQvXXCrTmowwV
Afa89mFxyE1PqvK6ksPfFDHNr7SZcO4H+zEWMqS7xcUeBVPwNGyy+BlvCOBY3GcO5utmpLxyPZXQ
HLW9mJXbVVZgYHXKer22k9hcch9dZqru0pPpMZgp10vZ7yr7xkuDyx6mYsVcqW71FyNp/kTIh2/y
hIph+f5a39IsaQKBVEyHLu0t/xgwJAtg2XNHgi04J3jd04g1LbwEheCY1XkigtqPJhU96zIOcld5
XF/58HLlDWQuA8lPftqkAUoTw7g77EfFu9cE9KEOT9G0Ptj33WIowJqYuLBMS7x8A8BouLBLthMw
IhtJsLDPnaCw+fsyFPCdZ/isKsdEf4YdOCjT08EThS1Bl+z4m/vugxjHPfwGCpALHXkPzB7BB8Xp
/cY6H79JrqfuwyFRoh40S2LNUCaQsggFZ8AaT7wgmI43KtrFEC1DMVFO7RlQS6Q27AN2JGCEefQ4
VxkEee1Hms3jerFwMMb+dDabWBGfVMv99Ab0KNwFBDrA0wOaJ7En2cT5LI6mVOFgTRrq/duKSGbR
J7Aj635PMZ76OOVpDRSlotfMEbg/FPW+uYbj7c9bFJ1rQHHct3LXQwTNlVePe6xRF4tiuJ0O3t3t
3uulJjbemymEXoixGyziHvViEPspF/q6nLjsTIt9q1vl0uGRQny34/l2Ou2WthrM5d1a8bKd6IG0
FtujHyLW8oMCmpJ8V230IyHxS7cf0Pt41r1EWxXPjgvTkSIjuh1V43/8U0E3WwkNyceI60t96/nB
wA8p0wj46TCH9HVzp0WSJV3eUGkm7RAKryT+fq7wp7CPwCdaRn9mBU77iaaD96yjeOiHZPUOhl34
BfexFXjdGJFbCQd4eEHQzKAmi1cjN1V68313RP/meekgeWzqrk7mOHw6rm/ChN2a9aRVL8niu+8Q
DF/vBSp6+pSgSwMYYBxyjyLe2872SedAYqhH2D/qlpAbC4kKDtWhftx4mV/bmb8aTIFJnEMG5kU+
Xwu2DKTg5/JiWIPzGYP2mCYg4z38T5YjNiZei5eAX0cmmRixXRGUZvcZI21rYpOabOpPZu8OGlbT
KEo+Nt3Cqsv5lE+QLdKBLrdmvVIv4yYsvn1qMU+nZRCC7QRm4vZbtD2cn7rGf72yyT7UWUPUxLii
53sSaf4OdA+mFJKdmTRxgVa/DhqzHajg0VqqegfFT9p7vqlo+hhR6iYJ7bnSxtzCGC1yCxDS5F++
uAvZ4VRzj4BHOcz4USZiKUAJ4Nt/cCgvn//NGZiiIncZx0dsaC56qFCNAKHDvqVPaL10MtPmEl5Z
ZVUFcb9PxSoOoeekyPMbmHl88Z6AhZusX6TmrgbOJc8WmZjyP3yowrykUJ3HpmNeFKxw+NWwJrDs
/rj5HVpnXXo4woCIvm4iTx0taGxtGOqZCsTkGnzBG8TEpfv1kA7q2dUfLWnqEUDUw3rrfQT+WR7E
zyiLn0zd31gEdBI8FF+tQjxdmZ5IjNuXdFK2CeHj3Z/sGOhlkn3h0BwZDDBAIA7Kpv7QoYhgo6uc
4HVaN20/UKAzimfwF85PZyk94/7Dj26LtAVQ2xjUovOPbtYfoUFdqcrW29IMbYufbxLnobh/Qfv3
Rtb0h2spj4zC5cxQ+MgACxLSBK1w/HnK75BO06soQ9UV+hbuaOD1p8A89LuORIui+5+3DuQOo9IP
2cTjdc3o3EsnltdZxk3lXYoXF3HYLQM8Ny5NTDDZ7pGC/G5fsnJ9JFxD+Y8YNV0muW1Nj0r5m1bT
bLJTXegwHEZOT0g5Ox4kDFGJ3/MT2K7LGopxwmCBrCs1Nzn6IA11c/N7Pgx46z2zqZQQjHh9Ybvm
mLlHjNQZpVuz7nzr0qWfFJ/FnKemeTsT2sPVTHFTWLozJJrZYfmOEyHy6xZbH/LFqlTln7LDVnoD
l3inUdzTW6RNpK9JVqs7DvEKkRb7ZrgTBnrVTMlTSVfYkSVjKecYUzarWThVBSfx63Vnii+rhVuR
YuzRuA3Azqo/tKx4tw24G6IcZb1s3oUp3bySMDt6qDRtKFtRgskFYnfHhsNl5fGGUl0whyD6hnlf
yX9wCLEy+ion3GuN8xtCMP2j1mNMV0hfPf5x9vbRo2TeDw5+k7ECJRjAM4/RUfQ+BlAZcQLnLTqF
CGNiz+5mBDKW7ZJ5TiNGD3qn9ef+wpnGGeoggLVYgTfAd6zG1FYWTqSSsxvOQCmrN0n5ELxK05fh
OB9CVhZ7EOa/tREV00+S2YDSt6sZ03CLRcvh6kVwIb/RK7G8SG/y+wLxWQLy13Jq0jiAjonTBoKo
1x09MkzILZa8pNmAJSny3L+WwxhuTY+iaJQ6+rHc8PMv5a8Z6/0zHEJPQKHHOfz9Vht/CR59ZYfu
xIGYaiQWw+zA8ha3ZjNSH4EUFHs6UvvYp2gWnQi41T2HxeeV2N3wmm6tbUUaKasitpFPIyV33ww/
wONuzIl6iyz34gNQItzjV4XhSQA9jbBmaxKCshDbqb9ugHjLDLtgXFcOBnBktqFKBWUrnFpojPdy
ugHgIilpQe8PcBFhvUmOtJCn7rOLw0r/ZI9HbKklHwjkTkaWfDI0mG2WoJcHqYZydURvrC3A1WBv
WXecdnApHMizgwpyogE+/w6yhVE+rBvINeEKPdCMo5Wca4pqQVlXIU19VzVWjBjc2gZDyt+cW2di
zowDQO7KGItZWV/lb5xDsvxeHHL9Z9keYtSm9hZ7S6UasygNyucWyXmRth/SbQAppCS+BwVG1f7B
lwYp1/VYsIK7AEmDFY6cUFXBySjzDoyaAmGzX96UT6Iwg8WFPiue6wcqSkigJ5i3E8Fhzp8Cxh/8
1PCYpzHyjJeiSghMppNOus3/ejNaYYmapTR8GKV4dqaOYkvuNKAlvLnOlmt5NIizdWWgvLV+aUWA
uSy6K7IUYGK/CsNOowy2FvWzuf2raR44sopPA46g0wE+sdsbpv0l139xLkZaKNXjVELz/Ke1Sa/q
si7NFYvdEx4BAUDNj6FVR3/UNiqhFDptVTbsNQG5LbnkXr/39uW8B9O+pENQELDGwo3hnIqQT3im
wcG8hkB9L0vc+4cx85mVqHAPt8IfQQAGEHW1NA+THxGFUaARGpvfzPku3c9al58M+A7h3HIRonfm
CAA+eysmBTW8/4Uw8wdggy1ubKa6WUAUNAKSQCMbx7v5vYGH1ciLHnwfiAnU2XdHwjz+Ycr6kGYJ
RHb3jBQ0KBaeTMWRrehF1OyPaiEMir030k93OkPIWoJD7DQsf7JqaKOBPC+toWfFf2LAq47h53A3
mW2xxfrrQRdTiK2BctOxtPsEQf2jMnaUporutnLUN0e2Ln/Gj4s6Wwb4LicA6Pimx+d3zPauuubw
kFF7FgsMQmAsrTWY52WdIxMpgUDImACY3C6iUj6zdghybKrTsm6b1VG/zq5qmnvC/NWv/jhsr3Dj
CKLqRMLQit5mdnj8UcbZ86vV9MrOHZIdiHMqJWiOKOzRfX7U2a+Di2ZZeRB2hG3rrPNSvVirf0UO
r1QQNt+fYVcC8hL1uEX6kEQIPifAXs25t2b1/sbHjHYUODLXfqjDJmDbjX5rSuc4DdBwi7Aev5SV
PXnlZvDBVb4XeGpksOBrCVjY/IusNAeLDZOUrte5WAU0XYSLUJ9gGjstAL1lXjtFq/ry3o625giM
Tf9FPGg27c1Liju3rI7+Kr1YolxbZgCkKgG2/mXZ6VrLoLIzqJJ5hWMujY6aPHvJuyJRpRm2qFq3
gEvFL47AsOwvIEJZvdjVwW2SLal/sE57n5vSj8UKuApx5SB/Gru2Pt0SbSDDbggF/Qiw2dN+vgR+
AzmgsZfx+/aDodud1tvLtcG1SiRQA0k/tow30RPxCI86vrSS0HZVuPOAIwPZrlJVMaaUBN+dvtS8
XzcpejGF+nyQ6Ph6t+rU3z/DXwjkv+tUvsX69EOY6Y9ZhyR85ZgZKeylmtNTlMfhcdGvo8TvuYGF
xTXf/0bGWTVmtaO4r3TNf4SMfWDFUd0qTxIr5K9b2+uQQcTvJB/IiCyL21x79UxA13EaUN2A4UhQ
5hcNRelsDBX1BiSmA9fTcYXKTfr8DYOtYoJmBdGwzE8qbKxWpfdQKyoe6o6Stp0ZwnZOrDxW1QdC
+oCRh3UxFsS7UsKUyIbdiryb6XFJvqHQiXKQEAgIgRWWA4WCMG+MYx5Nc0QOPIDj9y+MqTaABFyU
GG3RjE4FeoHP8n39KCSUIoBIHt+FLodvj1xdbGSKCDkBRBAPNegJ4F4l7P6n/iERPeOdWCS9CDNi
sBIdd3x4RDHsqTMQCoxwctANvfMhdieRKavzL0nHFByw/0P1fZhfa7d3hl7Ad5FZUTTP+Fjt16Np
dD5R4KCwC9kSjWPy3pblHWgnLRB6Jqkthq67SNFFXMMewS83cs63nvT3Dh/7TntRxG2hfRQb4OUV
+x6wwcjAHTho9T/On+ojSPcgxizdVdq2rV8DuelG0dp9DafduKuxfvbPriR4H4Gmk69sCIe/dSfN
pfUf471JuhZhjO9I1Ww5qIXfUSs+Q7AZtafSTfJ0dGn+6ygWtpNqYbZb2idZ1dO6f8UnegTxJqdI
zZCI0t5B4ENz6Sa+tZfwSCwrGpmPwH6UVaPv5OihN3VU6iQc+dE2A59k/2Lt+gQTnSHs+v5K2gyV
1EP4p4YkNj1h0GzxHalJ1tDAlr869YRvF6UBjFKq0BJAA7Zred6EcgDkQr70AAzCJqi/JJj2p//w
GXfwtBgrxYN7h6zgcvhoZiB9xN6u1V9t23rDUW175ecfRh7xSVCE8ko8mKdI4+6+xNfOnld1cUPH
USbPezAS4tRzJia5wzzqvGkpaWZgkhctpFRFXsfG2sH6mlj0HstQxpXbwHLxpN6uD1ntg5I/Qpy2
d7WF6cZuHPhv4t9jCzHAO4czPNCeDBGc6ENAWcPM1KJPr9AE3GhnDfJ1h0QMaRodqQzjHIgWzC3x
YQ3ASLEbjV3gP9q4y9aE3fMlNziwkbEhTmnVdPdgzMX9LkN0jzy9phCaLPUdVVELLQxFJ+SdLlb1
6h2C7J3CKvMP1FaPSdGG9cwhafjOQJkHY/S8ysujJmGrowNQlRrUzXs6DKIIEUlYK0XwF6YypEQD
gFtGL8P2+kXE8PNfkkqP4wUperOFwnEt+pCfi2s0kNcuvHxKpEc6oQOSpAkb1Xcm7t9NeITGfrhO
PUT8w/k6Le9s6++DH++LchYZsSOIOU9jCGleWjRocL4C61uNyF0RSUM1iW1sLNVnhJ2/YfBAFOnn
nhpQhOufFg6nnE7OlG/IS6r3MiMI9gaFqhG9QzPQLF2V7kI/j84/lYY8Ej4cEenqTXQE5PvLZtD9
rr8vUN7frI1RRg4NcLxjbr7+Nq6p/SDDEmv0SKeGG+J1f7zCaapQCYobYD8kINSGdSwVWP8n437i
aD8lumt3S/f2ADijG3N++B2bjyx04xRFnfvsAl0AfsO1seWQyjgabYiGYqiYxwv0Ydvw0moeBs+C
TnILo5Qf0YPJQi3Cs1xg6iAWPcOZkrE+CiwM+NQAbiy/2rYFGjwsh6AszkL3mhlhs7lbUEND6ZGv
y1nhZocTW7sSYeExbYFx3KPg3+AmJ4mOiiW5/p92jKoLL0rBtSvR9R/pd0GlLHbUZfN5AjbsE2CZ
v746S+OmGioXyBTc5JmKsYKl6XO3PROI4S0lPqL9TpiUlS8EAL4NIz2zo/+qDOlku3xgLY2WMOw3
F0BjdJ+BeUeTGJ3B5wInqSmW3lQZYlpDX9gVtG6TNsIHbckZqXOw9hpIV6Lve//NZFIbe8XTnOzr
1E/j3O/aGihqIaGLvVd9vE9kGMD2XqTTThbOBhVQ2GXK2JMfgixIfnCR0xMv9dcV9UyiGxYGw45L
bhkzA7qg+XR+zcs6c8ccWiW5eASSDrhqTXlPsrRQoNONBF2U0EDvk0oK22ewwPNoRRmZvD/tePqT
xGi+qzMUuFxA7M3UM/vi6r/fsEiQW+zn080f2xCfWF4ZRgwnDP3Wax8eTE+n3cT4A+3UZo4sxepl
sDGJufiKe69obMb+oAm1+EvtqiHUWQgClipY7/52YM2uCV5MB4OSsOuBI1EXD29W3DL6YCSHFh+l
CFJJAZ5eI8n3UZt4gPHneYkwTGsh4fD5rD025MywrBx1sk/NQZV/6LjKcMDqjtIoY88ycVTFufTv
UscnTu3+UmriE2YKL3Pe7vi4ErpPSKjjdi18jRZC8aOV3vchjp8AF3e2jqTifpneU1PEORs+Yzp1
XvYyx+Dvf+R8etJIZtYNl2LySqr2UONdQwlbeSRFZv5m6eM+ccHPa2UI3EgAWpoqmCf4TIH/uqaU
V1h4jvYXfXzCzzBGPgi7Vlp+xeXwhvO86foL2/kijf0ZOUgaEuwflX7q25PLRDW6JeCtn81EgPRg
u49rM70tyZA3WHYRMApc135P4AsDjh2LQ824w/O6bRUbrp4mxwceIFiIGJEKwdqGz3mOhcEQ0n/T
dBZ7CiFx+fnPLKzWwE+dpdz9GU3BsGQMmysZMDV7cDC6uGY0+iv2CKh3Ea+oyg26P7s/UiMYyz0W
0K9R2z+ONolb5kgPi/Hr8G5wyuFdGc2pTQVgEO/jpLKmkgHBQZFCQA3jyY34+o3XBM4ytE1gCNSY
AY2mT85nFv21N7EyAEMiFKC99cM4uEnduEcgD+LKJD9BADoehWm1aRQewqsgwwBkJMrC8sjJ7dfV
zUn/H5EezRk9uagwixsm+7e/Al9zyCWuuDTRUFFmsbex8gZbTYQJ0fGGfdyBJoX2tpLhfopub870
QV/Z/LEKqNwZrBWUcAZlfXO5ZWOKKkWsASD/xqEUC8+p8mNB2efKLWyo6E1Q6U53Hwby3g1v/AB8
wTomb5QPuti+UYjRVMset2XxNm4pvcEcCr1c57YhAENhuMUV8K7ebd/x8e2atankQ5TWmKtfySiW
caJEmsqpZogMFq74x9gAkoeEk5Ud8UG03jtkeK0e8jxjAgGqqJKiV9g+coTuG4ZjThgBDtZ/95Cq
d53RqYppWta6qjvvnicmB/ym273KcFPXHMV5aPHw7IKupQQk0EZVaoDOvCdPhN6QXyBbaSdwAaBE
KXwz0xGUNGGea3BfGWWvpvBPzP/JlDeL/5XOztPOIFJDvzcAimeRVLHrey9W/qqdI5ui21mYQfXd
wGGytDonz79EA7KYLU/Z/0jh/+mOgVyksAaKD0DqJ1GptEUu9O3nURMmsuvWSUOq/+ODmQLVnTmt
mXrXs19naSYAlf8gYLqXvSpgJOWRuVr1w8IvvKzQFH4wroDG+hHYwSp3+Q/q8zQj0M2s8MQL1fl1
sOgZ9L1UBdxrg0uC+kdAhRA1XjWGLspGYD+CnUX+GufhVoZPj+rLFe3IpfiMMP4ArU3Dwkh/5aCa
A5y6KdZTRY7snja9Am4TIrMh2xYxs7WhpWLAIOtPo9BYBDPv6vHMEeIrVOxungfSkYdm0xAA8d+a
Cd1YhW5nRCw4u3IwBN3DbLxcgGz4Ph1nYaYar29Wnlh9MeImZl4m0fFxdY6lNXzYJXo/8dmuzok/
mj2GVAQlz17d2qQFnA0EgxKp27pz6nXR7LvVeQSj82bKsptameVWsfkmM7i+JMPvAAHT02DF3u7P
QQWMGZQoBw8ij9i3rdPwoxo8itn408A4dFbklHz7yCdKBdsb4Bj69j2u69YOMcbo8cuK3w7Rv2+W
B+3v8ZyRB6zCFVXFICr2kRo+WyC028MYTyWWZnGsPBTrsyG8ACQfl0d4G71vl//0DEmFEwubQiEj
Y7mUPc7Y1tfZiF1NN2rx1iNfeXL+M48RKIYwBITljVzTzW4Vs9ty85oS7GcCjs9U2iPo7irSIajM
NRUXoxoLzqyVSyCvFwhAjz2M1mgWCUVYK1VQvSn/P53BS+MtTJ0nwIx7R6aYsOky12nLvodYpJkj
muCIr/HEz5aqvPP4N4CR8j2v3M2upbIQnI29eZQJ3DhGL0B/95i9nC2yeK7VHrAnvXtIKG/dOJM3
0oL+dMhe8gOP3CbozNQ1v82NcUfUSPxURgjhc0HhvJK78TwoSnY6bC7huogpGvt58kS8EmK33GwS
tcNIDAifI9v4EnYdSARq2o/Spycy6J25C2VW45DaolkxAv0+8SJs26yG2IqW2E22ah7Owq50F46X
azuOZv9YNtSO3U0Ta4doXj+XVrHlQgkTrm8El8R8DEIG0bbrTKWTpm/QylOfIaENWyfKymB1CdiU
29IVwUqc19q4BDk2PhlubPoMegXA6HZYgh9Yody5+DzrGB3xHKpQRDas92AtJR2D9XsxRawHfyuD
InR3ZRAoO+r4q7iy0pMfR6FSN1Zmt/e5KiueKjrKGJE6QIvgAX+FaQax9CVgYeWnUJ5ywg5cSe1r
ZPzjakqv0P+cdBtUY0h9hEMWyTz/rQ9nuFvoQlTt/DU6eDTlQWwpJGa5MUFnoXV65tGJpkN5OBaR
X3seBurtO+zweJw7kimBvW86jgeVwKV2vqtPuQHSQaUefWY/0VtxRIfKwb5zAsvI4Pomiev2VX9z
dgkUj6+C0CCuLBsDKj8IEuWnj8gcy+3xZuoke/V2i3wkB4rhY7zEdLXjcDLv6E+VDmpGd6SSu6Xm
4c4am1ErluLA5AyZwM7hUMVnK7BgvW37e2f+1rRfdC3wzdPeovlO52cIfFc4i/JkbmOGgkQjyM6m
xqBgdRATKwGAWYTz5eWs7M2VJXwQrU7SoiGjioxRKCnLlnDdkkDJjALoPPwd5vTANj6QWIuY1VdH
2wS03bRAyTpBm+boAA67H3cYLXiE2s2vIvlKYQeenL9pSbGdb6e3TCj1fO0oOcRW7KPiO/R/Pj5w
4pLAvLzuGA1PmgccYTlIMO0ngDZy8+k+kdeqAnefk1K5hGLTQ8dmYlRXRCIUWf1zr98nr907kxh0
7Ngon8bp+T2NLKIsSS/LLqR9mwsbI9P+kxqBBTZfq5sg1wvogRqTcReKTAItwC8yOq21mJ9VREt9
JAd+5uVwR0bWlph/BFyWl9X+ohN4mpdQAHbk6f912WxTgEDGXQevJ24TRZTz40hwYLxgeVc8S8uS
QiJBT8n/AtLacWihEbfgNB4RmiH96TqY3q6hntyzk/zluRLY/uVvAJET/Sllti8849xRjkOc8XRE
Wt30r/aT6CZqJs0O3EYDEpV3SkLylWKzpwvyZwmi6lZtjyhRdQ0bzcGyiYqIWoA/z2ZbVK7ATIgN
r/yi38pYRia6XJRHzR1IzAeZrTnh5/GCeVY8khUdkvkuqeWJXLkW8sCKsfwvhInsIzLOhauB08ca
79RF3hRczFm+Tkr2SD1EmQ9uRG34MhEsloJ+yReGRBNCHGb8qEN0m/GalkVrvsHa7Dvj/kiO/u0p
BeusFRd7pvaOQ/D4Y3ysBrutrygO4+oOUu+ypKFKewofF70MwcTj34XhhrVgAr3Q4B5yo6dFHO9i
lQvk0yLUe/LXhlEziYTVbCskmSXjEpENuZ4vmjT6kTroSbnYdCC3Ehxh8tVCYzS77ay31e41ks5A
HF9Fn+apkmGC3jKEL3VMUkHg3TC2dlEeSUif82zH5ohEALR3b8k0bqDfbtPN4PmX3eg8ikLcrWEj
kF54nEcEy2t6xUXxW4GKXBldAOaWQx1p6Z8yKe5Ij/Vi10dxj9piOC4ABThlwow8fsbL/d3hBxJc
EaGze4Y+ZgWlwsf1CoFcezyH8A8QOPxGbuHwOucAxQFzknNvLMf+hNbqw8f7qGwrjAp2BhUVfDfk
jmtoxvRh695rJcmrowChEPuhFwVWdkuIRL/+Km6LNSgsD6mg+rY2u6UmF6iOI321L5Rd6lR0Tm3o
rxElNd0BQcHiO+gSWF6E9H1oZQxDdwHWW1z5zM2WrwDqD3NTD2RFkC1Ct9eU+CzrSdYHkLGsIomQ
gffZ/mpgjrECXlhZH05aUS3AXdsBYvKhq9eWPNWD5LYnJbbgiPz2yYGbinCjB3JBtFS4x8TD+zcU
suGBWlm4GTI21/Xye07WzgZFPmFgRqDufx5W5FgHGKBWihgHNETEMHR3OkMjT6Y7RB6fq3qWugOd
ERuujYL4RJJdbJta0l5jjPXEc8BlcIgeC7aWfTyrr1Z6rlJFJhSc1/Iv5MKViXyaOrT9Mz1rE4R5
ood0olClj33q0SXb87joZaPFB5iDmzv9c/XsAUtC8UQjpav/LZZ+nNo33aXrWneRbDbx+Kkp8Pyz
Nk8XXvVphi9NAIoEjHjrY69tCSTRpvtfaXDjA9SCfKYR2EiAxqLMO1r08svUh6RvigXImcO0EL2y
dQ+az5yEgBbDREqTlIU2nN+vEtzlMrcZPSjNALIThkQdSlyAStDltF9xo0XCxQeDuCqWr7EEUZwB
jPWngisY8sc3wRmdy2XsqQspApgBGiD2oSqN/KUXSso5mXnQqA1lnyQFpj1hynZWfpCKXWhuSnlU
zRmXGNnKnl4Az1StqHZWcwlIvcLxUYVL3Sz6QGuExt+4fsV8CAVbiMNX7KJf0eDcL1zLfb71cQPF
I0HRYKlznEqDCpgGOxhSZaOgDgEuUW4hpSovPQFZe/sPC+Qv6M6hGOOg9i4UlXGPxaFx+UQfw2pN
J9XRo6WPZwnOYH3YIaNgWWibAmPFGt8D5GX0Qj9XV9MdoeDkZ7pGHB+FfPSj/tEvRg39GMyfdXJP
z1SoSLEVhdbTxeLBbU0LPcO4/QZAjbcwiwZq9N3fdQy9CJjHy6yaeGDfi1XLp2LCnafFeXJUBas7
dyxOkEaQaKyJG0rClo0bCmQ3l6/hXVAGeboQJd4HQv8eW/95aq2LzfkbyZc6n+KJRLzTneUGj0cO
Kw+5h8rwKPZCDae/RWqAbRTy6MsheNNWf03GX1Lgn8mcHfsm7A0pqjYsxQWqhB71IAG/IfxvK71/
iSqRIKUbMntVKZXV5qgdLGn4Cs1Or6hr/2ndfst2/SItstD/QKKZnvpuCNnxxEXQ+8hJVzuEPYPr
SpeSTNSlqH8hajjXy3t5URqtLO9mZMsYU4kzuRwYE51Kq8ty5OGP+0SiBY2towOF1p/Sf9115hXv
EBe6jiDraVhAPZ4HpfsrHvUs+MeHFmwfG1aAqpsRqGAUyHbcl+D9nu4QqNrygAdLrl1F543gKraR
5UlWpdDUOLyl7LGgQDs4Dg6gfGtycTsb75GP/PSxeE8r20A3rNkT0tt482uWnv7wSSaI0gWOMGhV
OkZFqLXbeT4OIylHiVDTD6EpMBN3SneJp1QmLR5Xf7bSYPve6/NPcIcn8okHRc8SSlyMuK143q7F
vSqPCzTnK98/1aqfjE5j+AhASr2HWlNCfw2SPBWVtZJYVaFxuBq4wfTafD+cHATFAQp92ZdhyIRP
SMlmPHZzbf25Wkr/6b3JRhtm4pPgRo9d7sSRkjDQbktVjYWWUqNvP52wxrZesK99mzfYnsJ8hfsv
Y2myJOEbJSQ5mzWOhPOYGE/yZyn/jlGE0RGQgQcv7qEgs68HO2KSG8np21EYPE6XKieUa2RCXh8p
fs5zdAMtGQhuP2NPB7iTRnSwomkj8WGYPmGqKwBFxGe2FW/4jLRzzBl5rzJQZwlGvm4VBS2F6DVQ
BlBsgM0Q9yw+Wz4n+sToumPXy32X1YOtjWXUN74X9URj5UKdrFY3OsSaVJsyGaEuYTe+mgzdTMXH
KD0OIJwkW/nZ0u5jjpD6d8zvCc7noy026ItQH3f3ZKUiqaS+K9uKqw13Xv5vuSqT4u/rJ9KCpizn
chdoRWB/qPpIJCHcbqGbUkV8vD04Q8U2TjctO0DiRXX7vz65VYEo6d7Dso8coyZjskaItxYVswWS
7rqzArrG3sTNENdhBoJECh+2zIxRf1ktRmySqgWToVno2eb++qxO7xpDVWIZEnaBvj2DNpPiK5tC
H7yXN3FgizxU+IP2SINGpXVkgUMIP7JQo9R520yhD6vI44lMESM90sPNG8vTBUQTKr4BT+KbXp9I
mjO9CZm3z33WS3p0EL5ufrDQphAsy+c/T9sdtU3EuMHdOY6vZC1JTQ6nTS8lrBDbm5pbycd/jp4Z
96/kNeTBWVk5Ol/ZtseFeq2nOh7KxSP904DWfFfAKuGBocIgYXIRRHqjsUNtlSMmdBK3IQUXRya8
Xk6woKRFMU1Cnp3Vhecu3vr20wEOCZ6obr8JN4EMZQOvYKTnjmsRUWmAlOHRdb6IZkCqhzxUTZE6
sLym/dhIkXNXOPel37iqYVZPjPJKs+RbIhFTJ4S7uKyhUPBPYxFtLPjiUpOumNp2yovFHRJ/AO+F
YHZWqXHZjJExEn6Yni7Pg4gpu/LNS/nSzNhqaVOY4i9zhlZa9k7zjVGRBzLJnlH5TO1ck1smhDob
73nrwcvC+/8lyAnf68JoBi652Ekw+8FzSL4a0Kq0PiERsbyk47rXf0ysB45c9aoNbGaPAmMIoia6
aTSo7vm0e3bhIBn3RDZOwfxvwxCbND0pFvDBM7zaamdHX/y1Uz0SReuVK6auBaxtsX6Xd8TqgRFp
Sb66AW0/musxqSNqSClnHqPqN99woEG68XKvd+4fSht+vnHB0zxQU0nEda8fz9iWjodAvIcPrQry
DrtN7FvHU5UaJtYV94b4u+UHiy+mAPcSdITrH+RTHV0zqXu8H8bIp66BwnskEMwOqeP96sV96j5h
aGMUlSxkyFkxmHfRNgEXlh15ok4w5xvWY68SOll/ZCyw1UcWortR9RhhvmRp3WAZdUiuvhGEM+5p
w2JFSzupb8wPB/C118SzOtiJ2Ex2bxAGyDbnY6vLPDO0ALdWnFCB9bN378foma35dIZbDe8XdBAQ
PyPs5AuUCQEG0++LLH0WoXXYEZtrIMSl47WsNfC0k9SNMet0FLCZW8aBfi+bViLjYVjB9Er5xPzN
rB4SCMstPiXFOGfM28QnToXb+Pkmlvz/GjTDCV/o86PGTYKnhuzzkrb18AwNImw3p9MfmgZY05yK
ww9fk6xQDJkK0g9tF+sBMOfAnPIDeA4oOh5LmXP/gYza7/l0wQg2jjJ9+gh1fvesn+sq+Ubgow4K
kW9hJeym+N2qvBRcCNzjY/EMrDVGd0t27FXBD8j9SA3wR9AQbWds0v7Jt/CiulfzhAauH267lsw7
SMxlVZkG8zhPM/9qidvCqLlUPYlQjneC4Ix/6FCu1TrySQuBrPBKrN7XZNJjZOc4yrs3nEpn6Sy4
+XVvzDbK3dFJh0+gqILDoeDdXTx8lNXQd0DjXLXNpOQZ65lKa89UEaCtrv/mOk+cvPT2j61Uz/H8
v00C1Y5WCTImlXsdSv50ifximHYOiW0gep1/quvqTk67JEbD4C99rKFUcZPpqIEVg+jBeAj9NPgZ
DZUaTStRWqUCTcscAVYGInGSpy7EUf7hAA4O6E90Ba14tvbIIm6xwWrcVe/eId2gqgYm+ZkdPOCB
bTi1FAbX/yFaGo9QF6itXaKbYVviPC1AkpuZbwubQGNGFsAHl89pelh09gSY3Bk2DIUjBUD1TZcq
h8pMQ0j16xWck4oL3/7nWvdoDLhDwSW8gCtdujDiqaoKxTBtbMXSlcZ2AtLygC5S1k6u8ca3RKCv
XHPVhB9+tGg6iL6Gwovh48Jb6F9+BPDf8rbEonWdPsY15LdbTYz6xotR6VU+BDdabBnOVthjjd4m
iMZZXfGpzKVy5vcumR3mf9Mubu8sR/PMw5WM3b2QEIU1VMDjgaKmmJMB5HGQFoS+++WbdWEhY/Sz
UYtFNB7THPgU3RrtfKA+eR7FzTZq5qF7weNncyvvewxCk0LVxQiKsEPhEJMHTC+ptMrRYfetSajj
Gn+Q7bD+wVEf1KEa4bIzYD+1ntcFecWJgOY/8ZrUBKuaLHqIQueeVRgYtOhTIC5IfUJGVFT08Tmz
p6Uj+tPbFljLWuSICiZGeYMIZDHWW4vRTsnqILzQAon1Fsm2IsTsxP91kW9R+8Jru2meJg49wMTE
DuUpCXLSoX1SlYqjfUuqaDXWCl8H5QuE0dU3W5Zk8VWtV7g9BNGPpjh9irau6ZmBRtXi4IXzDCFx
T6DcmLO9JoM5EjDrv8qpaPfUK8cTCUVM+NRntyxek9bKghhNw8WRubLGfyDOa596Aj/epQTfgcfC
4L05WOqmAXO4mCfecnJhtwc4eSadTUla08PBsTNdZq/NlfcjhcTicFw8kTX91EudBnLBLMr20eIL
qBCzoKmsdh9KSkCheAUW9ecgi89yinpcsQJNCww9jYGmjFNjVDxeH0JVKfTxBXwx/nb54TAsF/QW
SVKG2fuOTK1VG9I3k6cXnGoDRFu+y45CgZD0F9irsDlK2AHYbEmwlhLcZSNJLm0MdGYFPYd5bzpf
3ny1xZCh8MgpxmCQ8813oF1JG1xHBYAGIhwwNGlV8Djwkduq57+pGoiPNMxBtAFn5mTuvv7oF683
gFlPZUXbJ5sSavgqxKof83iBwBi/TBi4o6UTYaW1YZBlzFLm7+72shySrpfJvLg3Aqf1dpxWFHWO
Jgeb/SE/Xk4PcqsofhK+VAMbImNn3xPprv/Vk1fQy7g0zbjCU+94GNL646V9hpeLVBdc4VillaQd
ETczU7K2CY7ypN20f0zQ3e7e72JOXE5zgrdRCuicwKwSc9Og72PbL+oKYEUcIpsPOrXN76UF8Yt4
FaNpTW7iPw4tDAanrxswK5lIwOJWo4JShXQkANvliYZHx7RrZ3MBT3Al1I65kc0msvr8zuElxetK
7doTyynBpwjQI9pwDGtYx0CpM7VRk21w8ll00T0dbC6ot3Zqxj0jl2pWucsoMZoYbG7kq0moun+V
UOUEnxt4I8DxD7Iy1nra8AFLppSSsHTbVUJXWohxeeEWn+HXsbDw1S0RzOfN5PJNN6inZxHtdSGK
JfvWtBBPJscD9h/448Z4CAlUFGptvIkCzYmC9uuxVbL9etVPavALgbX4b2PatQ9bl+Wb1YhmgHAe
QMRVqlVfOHqtjQfsCbTF2Z9uGEIS31Uegfuyl+EGbRsxGR2nw2uNtxlp3b9C3RfqSMgkWXFbzK7Q
xPx/hnvWu/eQoEMaxC4GHi2IO929TTMklKoYThv8rK4mZ0CugDLhNb+B9RIXT1UWgGB3iAeZJeS9
vN7lTGlndY/5gsffmF6LpzT3+Ca4eKeyFP8wvWplNzSlRAv0XLzXGkBAVrWv/LZ7pUG4bgqnuku+
JBC71kTKgpYUPBY3rl89whCRXbJqJF4br5LGHhDfAho/OYCzHCwQyuKXOGmo2C+mttRfNoSCNWjg
u4LfBY46icjTmMvLJZIO22dTpgv9Qnhjpn95480au1D0rZQD6fvQaM7H+gpwaHqoWRqJntxP8mIM
yXoW5NkyXNfDA7813BPXBhQ2eOvhItAQWwyXSiumJ6ILN7hgc436bgCTyHkcYmRFGGNtkF2jCs4z
PVMKv7ifydCnCSElfQh+gb6SRhiNPVovuzofd1RJuYml+t5ue3JBGz9oOgBVmz3bxRjfpBwdj6k8
kFk8lSHYfb+F+dceacc/Jk2B7N8MjRvhTzh4PQ4jdasH3DCs0l/2EXc3GsNSbKlonF0dDT4jvk6Z
8O/QQa9nVEjRK2DPRAhx45+8SioXAJsSk9BRYbbfMOqImZetK2cGcyr4IrCC+Qm7JzIYvn2Qpw58
sxKHEb89R5f3mPCfjFdKFVYAhy9LCNW2S2ZEFmHTm50i5mxUO8pLOkLNpMahOlyLDqF3bMesx6uE
uLdYmlczrlRWcugcXJEplC9lbpZKOXNZiLrOO/GDxyONkp6RY0dthSwiX0GIGMDzVW84UkKKwmfp
PUhCnZSQYrAssnPcDR51gyNkf4kkNe1p2H2RmGGsPy1hV/qk7eRFC+vFuaFvnLu20A8PHdKIMm/b
xu+DAOXH4jklKpO8SO49gd88aguIJZX3nCCLWe7Avilz0lgJHPttjHsgYaXOvxeBmIFFSHYQ8nrX
ChvEZhNZ2YGySpvKycIedLGrr5zXLatJl17smsuq1ZC1W1vzqs+AIFXqB3DTiOayN08KQO016zBp
SDDWv+hWaDao8avoxl5w1NA8zsyK6rXbh685SSzj5q9kN5T3D/uKWkTR2TjYgwDtEt6FvY0JiZkn
DHkIYKXbNCiurqAEm0jMP3IguZjE2Sa4cJHcGkuroOMoV7QoPKtE4/g6+npySxYYO7u7odu3Pcl1
x1vPTOzi07lMHLW2S8XqZwAxQSVl9lczdk6w7px8SPN31tpXwxn08/ZyCY/SMbaOXhyZwGjPNnxK
g0M5FLsiGs4q0pxoh6ZsTJpBKJlnpJReo0sx8/uGFlcmtCxL9OodK2rc+1QaftpbcQ2D90z7bDRO
1sonjKHd3qzeFj0M9imKqaKeGjaOpXwuKMci3x3OxCZIl3IAFHpK8hiSVzokv0JYDN4eSYrpsFDd
HJwwJMDEK5zHjC5sXIUnoDngmgj/7+mYqI3FukOQQaMQaJDvYuR6MIBNNCws2VQb1J07/ykmuFTk
loLgus/Bc2yoDlI8ycfczZRst02b0cbkHEjEXY7E7qF9lmU+pyZOGnZlKv9flH8w8DpHPiqWXtTy
IBORLgoumyw7kFFx5tSi2tl6T1vqaBmS+Dl0TnxLSsDJqYS5uh8TU1KhDeLUjoMO1GxoogL36e56
24anw7XrYqyfwCVSB1Et+qP2x+x07eEgT7Z/RlwOYE6lJFfkmMPOl7p8/sJgtZSBI+/n0zcB7yOL
FJUq8se5boxziTonPm2HkQqGpJT6XnxlEu8uAahXK4B0LdaPH9OQOFyqe80VAYlGWztHv0Uko8oB
FwFgsNZsj3gnFQ3SeyiXUOCIDPEDd/EUv06FvvgLLzgm8w5mctsfbCzyza/8zYnXVfk0xuGr9v9Q
Q6NaIpdQZu6ym11e/ghsQ4m9uhRCyy9PkzWMalROhZtwGrCwn4tJc6UizqySMPWtouMcPXW48ZIk
0msrgeS2XN+yRdyer3xW8OktDAKmfmXpOOfB3UlcOz2PB8klLYsfdaqfs0KfLZKEcKsHwqq8pQpY
EZ5S3Z3WQ0LoIR+FQrOVVdAVCHMoBdPNpA9Y94MPr0HBguEV+0AyscF1tLBvW3S+FrK0RRzo5NI8
pFc7YK5R4gAQfYI/1sf2z5DP0oj7nQwwlF92FWubu12msBJ/A1COhJ9rA9MkX1mc6hLuIbk3kj1N
KLf74aa6RrNJFqwWM+y9WycUg3tZUcgdKbQaY/KjDJP6KMetxh29uqDkU3MkNp27VvCkR5sWNBgM
GcmHB+YnNcSC7hetWK+OuHRk+/klCfHq9clwZ28J6LGsZjKWVoBHLxMTKVBQGMnt9ooIzAiLcsd1
gLm3jWcRVRFDTg3zft4FfMFu65ErG+AHAP5VsVXXHEbdePOkg4KByn8sOm3oKiCKN1UKkRkJyCU8
6Gq6WPX03BPyn9hOBMHO0Dt/B9JzTFi3ocaJIFWj6XJRgS+BqzO6z5aj4z88AYnxZr1tKCzAkGeJ
2zcIncYd2S5bQIdjEZVEG4+bMlrRwNLx45XxwYhr27Kj9BpHOCW3wQhKW8toEq4zUbTOLMTDl+lf
DDCy9whsweZFsnYmXdfhiZ3RcXswwNBrNlk6einR//fIv385zaODkjauBM8+sR5IYZHRA034n2Fn
Ff+2tbUecuR6kzfQzu5q5hQWqW3RKwaA2pokWKBtLjQ73mglie3eZ8V87NUOwJy6dXvXa0W277Bg
XGLDdWtPcI3kztCMIf2DT1/3KFiu7UcU6lgbrsX9OVsBykSovOm3JXMIsvcIS7YTcFRIxBhIrYi3
IUN3quKAX5moKh9DL9ugoggPjTtH12ILDAizKAWOH3rxmAmVBFfY14gJCo3chpNpmBBYsD5zWoGG
ILzEZspaVL8MQmBITNCR/+W3bQKKAOd2OEHyjURyJtwVBooanj+rgkRP45Av1mGklkL+suGea9UN
AX5N/MJgU0GyLMSbYb7Fgr6TWGropZa986pi4vlb3KrD7lS/DMd0GgDHOdBz14jCrmh17uZIkcEh
QpTic63t26QsADNe5DvxYqAPOXpDUyDsb0VW2GBkvz11Kg2UqTITOLYWiS7j+zrwIQJ6pbKeEY6d
N/oFn0MG5kmU1vYEQQYuobiGYKJUo2japR4tlL77gZSBj6xyCPG7Lc3ubCfGP2H+kXVfkLyVeomU
o1+/w7/O1R7UkEoD6iN8TEYSQIjmRuLOew5iYT7lCMIHqT61GUbtHuJsGJoPEfb3GSMcgmLThQCM
etwJwQ9qTbWhIY+1kOK553SAOLnI6vI4XI3jCXNBHudreLDQHhif1DE7NNl4nw3BXttSTVscwPdD
4SRvNNueje6dyknogbCz7+c03ZHcW4HvmNorSN+e+8rAj+FEVfywTE7plab56zZRck3bTMoXHFZR
KXx10PpoXbDid+sLA83fg/yXM1fkI8qU5Uo0BJ6tnEVGRJXmDamrcJ7ltrjNV6K3VQnM/34aZxts
JbKqQY1XirKa1wrubn3tIineVt0rOEEvmTV9Gngku5nlhnPn/2788GtWh8jHsjd+v6Ts9btFJ757
VdrabC/eiYSIux4jqQPUV5wrrwTDMnfoTOxxJHrIjkzFHVarbDjnlk7NkEa4/bNtmM8f8pyCUIsP
3HvdQhCEFTGvguwnBBRn1kvtt+y8Pk0tY2BhR/bH6CfBEcu7mQjw1yfZxbkytlhN8Pj4Zrr/58ZV
dI0RwT1KTO/0U/ispw+YvBAGlBcGMeMxHHnNDt9wjBBYE4VM32h3zH7HMnKXam5zU1R51fgMnnVH
apsb5D0IV/n+sQmzkT9S+RvgToDQRgaMBUElLEpAPYPyfOSzfLhkOnsqkl1el2NyCw2aqmtWQV61
MuSLP3KKdwseyOm3H2QjxoisYFGZ7gSP63nLZgRhuXmFUBkh+TjeZUlQfPceATtJhIAOJbFMY84V
IWMwqAgM40h6kHsq9owoEztv6bpvDUMjc6qRtxvJ2yQUktf/DqlWibpQ0SyBT2IU0CaJtEolJ4qv
+YRO9JTiKX465t+uOHe4ma5LBHKNck+pNck3B8UKz8PJYvSqn4w7BeQc7cAAa3hpHEOo/FRB0B3j
Ckgx7NUd8v+Yqo+JjQNpcEqnVVUFAQQ0NYGjbdH5l9q5jlSabApRBNZBvgvAIRrbZzFZ1bPZ0i7C
k0QzTx881UAhZYajAFXh6d2CA59aqkYbCAfik6K42YkPfCL/eSdMucy/ECU1cOoulB64oYxelvx1
Ub0ZpX3NdnH2v9xxh7xjI20sFxXYlM15dkF0564uPymjBIg0qKjaQi7R/1bXACVprqAhuP76cQr6
pCsAxQA29TBh3SGYYLfqg3V16NST1OmHUEEs/t+y3uufpF8EIGbGwJ11S7mOkFZ4WDhB1wezCYKE
lO1nNSEZzJYuYu27tvUq7Xw/edUttkT73V5v3VmlhFo9THMD6DKY+HCtVOCBls3pzyRK1A5i7CBs
DhUZlIvm1DzOZbHYrUaG2FZwIqVjAquoWqwuFLN0hd5XAsC7cAKujLXoD0q9KPzXcdavgbIRowb7
/AKcuijnQJNQZP6/T4SGjYbuz1rvqtxdnxwXKDJtP8hxf65dR1PWxmgaC1zsv3KNFMweM6fIytTp
H/VIu0WiOc6HgXtADkj6WQLuRlQzoA7G6HbkYrnp0ZHwK76yCTqUTpQwUOb5TezO2dLc4G+/9RPV
nrqlWONuTrkqcEaYKNjTLXXGhaxc/JQXAjrJzQnnjG3UlVXX922CG/iTA7r7EPrs/XwBBA0scMCh
73u2r1A66PZlk1MTmRB642X2D+367qeg/Y8BKudQZwiNDNv1GSqWcnAQ0s+nyjNKk+DsXMAp+Ezn
ciOecB77qcB8GjOLeQvJWC7bd9HqpxGFFZmR3qXHi2mwxFFPzIo+kvADjjPa2csxoXUKhgDpQ/5N
yxzfU1jDpOYEQhDBrKI4WkNvne66uS0BqB/4MKzWaryU7MzQe73R4L/zpwlk74vm7EdRHzosRAPs
bwfWwyJ65DbRjLL5l5d7I6B7h78djp+PYPW5+03Dmjy4ZTXURPVnZjnATqx66jgV8t26LNOC2H7N
p7BxnojQahiqoWa16dF0MJ8QkRTNSMppuXJESesYOlK5zkrHMOLC/4+rhRxkfApl2T+eF54KKM6b
Mr0TXGi3mUdZSYooDKjsWYUvOuEbYQyY5yoQjFr6nyWOS7knbE6ADlfDCCTayI/QGh0kPVPWKjhq
7JLo0B4you52Br9LbAcKbRu0gSnwxEeHsaHsOUPDBv4rza6OAoWd+K1w1FLTqLAgXCs/JKE4f/I5
jFZlQZMnL5J479sMh9tLTCf2QX7h6V/zwWO5VJhbxI2Ugn/333jf+eVedK+tbec+N7k1Cdrgx1wG
EGUg1Qfowkn6AINI9gue7MqVz7HjkSdzP+t3ti0QVHNX93NowiCi7dbum0d/pule6mBkm42gEnps
I3mO/SHOmmX2LV6MYIhMToZVo5IVcBrvzLFApm9+9ytgKRfZD3mgfroenf2L0Aw5UEC6LjsTrbcz
VS0gJ3IB75+0xtgS18H/B6NP4ZgOEKLiMvC41MQ7CvEtwNiPZet8SZt+AjnxUYC5m4qjcBfdscEN
QdT3C+/vR5Ub4nY1aR8pZK3ejQsg7UqdiR9pYTUpJkuqqB5qkqv2vMbJaq5CZRspW6pA1eZ7g1q8
UJDHkeCh6rkIqTfYEphiK+suDJQ2pI04DkzVX+Pk4riupv2Fa8zOWrkBARD32NkaRSTTEJZsAek2
004ncitBbTWvk4GkEb6wa+LDVV6dLYNcsSz2HtOLF0CNCSn3eyxwdLhz/gD6s8lHXAvC+Vvi/n8H
9m+KWZMvQV7uXPmmRh8UGuby2V3bBP4o2v/iQXoUt25ycwJbuWiwU+MpeqPUuAK4KBcQDuymbe1T
4kqfNAAxw/wyD0YTeQgyNoYMBu2Y2HR1A3B5U91tzGumP7k7oewGk/mm72Cduu1tHv+ovrKdlTyQ
fBDuLNqwb+ujSOPe8ktilljQp6aTbJ6DDpBaJwxy10FNISvJElOLxj02tXuzDhYXKY82TL/gu7of
TcH7goqpqC10/yidm8mc5qWhdcr7jzbtRePvG2/6NdJ9iD57iwK2T9bJbkiXrkoMiSuapUAeW9+x
tM42Ju9WhsZ0KFV3EN8lUYYpRBixWj1PFvWrTgcSPxPpSjpiJ75CDoLwEUZiJuOnIAbicwDwehnX
ryGYCvLQZRPJFtLaYi9OOyi4es+Lvr3u4r4r2ZutxRXiKucBKLZ2cWI9Q6WFM6zlXBOfGiXGsGkz
0VxtbExv54aIOEftOU2hpeR/XUKtW/nk6rf25dvkmj12wvBRcQ78gyS0nYSTWp9cSMs19Fc6lLC8
PsUomAKS3wl1W7MOGLFbA34yVODM2R2KD2FOi4bQJ8iqBPeRZitzzbhdvdUlC111Kv3fyQHtk2kz
6ftnlqEzzX3gR3Kj5R/zNqgJRPWnU7qT2taT/TohPnzMz7078M/bTRSwkR4Xh0azsJxKdh/6g3QR
gDbgbS4T+m6OVkoZpbLbF04Qru9IOlpB9mWLKDZeoRUpKo1HGIHV/Rtu7v4AcYRAMSUf6B+IKvNk
+GIzETUuNpda+ttzv3BFTExjNMxR0CKkxk0C18ISh4jMgdbL7m0FnlbnYg1ge0HDBLVmrLQCYYg1
O+ybU40ntoaj3+s+KnpKFSKhgJ15oBOdFGqSTIEXrDH0N4BT5YDlP1xTR9OsT4+kV+quncpekJfM
SmTS1jSOmXrPy5WMkqGAVJG2z4Uej9RInwQ7SJ3eld06RqGGeoBK/99NcXhZrJQrwFAdN4UCacS3
a1V7FhnewWUEUbneUMKq12GMYOXIghvAVs9qM418UDN2CDL1g9eR6Zqg+zQR4HGEQb84k3PlBy2H
751rXNNhi5v3FeBZtXcOY0Ctf+W6c3cftlrtXB+E5Q1KI6Jj7FMlkaesU1VPS8fJdB6LjF+Rr3CK
Hu6V72iOHFnLBHKPG/dr7d7DZbh4ETae2z9/2zLBvaXPVtJ/zISRK6L3rhuB1vb4IfFo/i2CxK9i
MHpohDx9iUy9qZe0XfGcqLgajgDg1OlNhpIE1B2KWXDnQPQHQNkIekZcLhigJqbz3FZH7JMp37G7
jp1bciwcoAYC8zT1OrQCnDA8M7MV6wUK3mThK+sJS8WzDxlES8zKBQfFBCWnqU+Yj+k8zTPZpG8k
o4ALfFqeHHwNfeDu44PJ4YBdUP1bpGUlDUwQhUMWCdqTs1/0qtrNqCBaoUF5WntVT8jI/JBsIaQU
+npOkPF00w93k1B1ykX9dHca5OO68F5w+RmwbyZUKovrfq17ssMK6SApVsceCnT/xfDMtU01/dXV
GGug8l3Jrq+I462/b4+YuPV51YIeguwdqvN0mV6vImwif+RJ+2mo8TBh540dDkZTf3V220R4AcPZ
uUxl7IJWwRStd11yEWsOftVJ//EeM+ZaYjpMsq0Yn3g/6BvhTggiIATgwcM0SmgXMImIug721wUL
ouBTY0CRFSOxPijh88xYT0OEl4rRKSQ5N/HM3fpa3tVt54pF7iMGPJaB4vm3SSHUJYrb4tZKJTLy
5K3vEwJQd5HoYCMK8XpBkL2F4P0rk2VMvbkrSPjapagt7aFk3SU0yqMV2g7ypYrOCKgeFHLdm6xz
AjLImiODgN6ljZqFGOkbEbxl8eq+wal+ENTSK3YEzPLWTWg0yYzbQw6aIp37pF4RD/ZmnuBpnVh7
f7ABk2cmv6Hw7STV8RFvVv5KgpQPwWWJo2bJucHgoxQn0wCjEpLqWQyYPKFl8S6n1TXe7ZXq/oFY
WqaHSKFvEoCRBUodu/60mD+nZb5lN4vBkfn9U+2bASTBFVJhO1P4EoxLek93t+u8ftLj/pt1MqbJ
ZM5uKh/s4elhe/qLeMjGPzKzDMDKiksWUtQX89KKGF6NSeOmLZaxORWucIzzOtNUhA6NXrywEJvv
t0OGygyai0kr+xG/TCVHOwSTgWzANJJGabpQL1aHBKc6sZqN89TMc2mFIfOtfj0500PHf0AeLlql
AvopsHuYi72dkEC+zB5w9McExkZwY/O29N0Nly3avg7NqrV6DAsesi7I83hzAzR0LUcxt1NUkakx
wTATqEh2nbt+sVSJX+KwYzvaIzxCOI3pFDcvx2UGXpMkh28OGkuAMr3S/EVwCTcVeAX5qYmt/Ak8
4o9Cl+WxxA7SGItRpDDU4hPb9wQ+7fW+o4w17r3K5ZyPUAXlCZwXhRwJX9R1yweW28a6ak3Lnzzk
G5hhC/DY/xsuRGwUfUTaf59CrB78D5rflzNgWx/LxpP98uWW+7RBc/wIzsrxzY0I0AZmQgla5/08
odCGmrsEMPOmDSoNNijoZ/I1otVIVE3Zo9FsxWaY4I00LRUkufI4KTJR4C9ZoDJHVAfo02WvPJKQ
FQCIzjswcbycfFfMefxd6S3oKgvZZX3JzGxZqj04NU0Cmgv7KQ+a5yNWb88OnZNcd8UhBmqBVdII
aSEyJXzrvX/d+/NPZ8m0WYXm3ErWvqMcqGoLziwu3zg+FRzyTqe6uc8KTMFHnjyffBnmBMPvba5E
Cn/F1ghhB3d5bA9rBgf32OlBiNHWqhP/5+vQP7BNmkErs60S4emYhsQLzBAdoE4SpFEcQdbSyzr3
QmzZoUUrl0DFxmRbNy3UmWSmhnOW5qIsQ2hHN4L9LHM3ysNkFj6qT3NgSsBcAlE/FFgu5+63Z27G
cddfYC4xLRM6v+mQR2l7GZexjOgKXbX1wAIoZaLiF7sQk/8vCERqIANcNFa/8YuZEXXf3rJKD4+N
K1yU79ob+p0Wt2/nBc3bZ2p56P6L16usGqDaKr+foGu9CNMO9hEcrb61+qlDEtNRZG7D1XGcTCZr
VpOBnahmbeeimeTS0oSjEK9/LjQex2A+RlYuDIDf92lc4HpDNojCZ1DzNh67ouDf0k4A6kyzcc6p
Whxb01k7cYaEJm16chmMt9oGTWfjI1goKg8xYUTVYaarTPNOiOYi8L7K5macSL7PWY+mYHQcfE55
m/cQBF+bGWeLxuWUq+3850ULCwbuZl2Ej+OOOOQbjtozH40o7BJLzAb+7dMlKTddeHsQ8GNspwlL
4B+zUDczUBirF/Z7JMCBeepbyl2sO4ojtL+v3L3q8v3GtHCwIbhF2A90VVEjsXfiBG4iYO/lpveg
DjYay2Oq3qnGYhPS5fowJQb+KXw6glZ5wKEBUWzIqbOpJ9IlNcvrVcOMBJqexkqNTU0yUV73uApZ
guDodZHZWPyoUycec6DEfAxDsvQMjQ7OkPwfPwClUPl6+eGQyO9wgJTvMA5N5FMO4deyT+B1sFLV
0oX8vLIWsnTng0zqk7ZZ192J+86hFI09xVrkfEry1M3W12AgrIUTaf00fHbsZFulYzwgdL/pL/Ro
YQGABZ2iUL0IR3bjp2ccLSfDctPxe5lVd2SgbOy9Z/MARvJUSolH3+UP9KWsLanvVQakdW0tPKWb
KPqx8z1DjGgwLzZ6yKsIrLuqhlChOH86ZnimA9uRlRi57h3TfPoenP79SAG05y5o0DbGCcdeIJqQ
EeDsIN80fRkpoTdUSS1xDkneXRA1N+W2hsdPh3qtiyM4Q3NnAWArPTWbZXRnXnTbuuBIfqi1/t5r
USt8DXmzJqXtkLNXPxWBgrNaB4GROTBN/lRHk+pxQ612axRZpZjfc5eWI/5psnz4R8z7Yoe2YWMP
GV43i6O36UXBDSmATFP5XWQZKbL1bKOd30nc+0PaNtCaKyif2nC5+jzxJeUDFKDbEZBXJ4Q/jfMB
zE8BuZosH4Nzze9aBZRzHoHMPM4rUiWJ+kqD5mNDNLf5aEolxv1KI/MgeX8rKbyEZpuIHXibI4Oh
52mvqlGrd/rffm4i94uT2hhkanrH7ZGWIyE42LYFb1YUpkBAIFwQKKzcknmLbWcrSuzqnno3ze6G
+NHOqvdhqFxuHSOHeXZjqttRiFtkKe9KcdKjXd6iX5LWVchUwxuaGVCTMg0AjZvlCOYNiznMHHHt
Tf8dkQUoHP/+KwrQ38lMb3sYiP57jo0yJTSwR1Ua5JfUyCoY+spgukE4KEYUAHfVb9KbU9prM7Pi
nacwAxw6LLWpLIOK/xRmGSzcPQkX/kPCUz+y2JG7LvMMgZ3EIjyWiFAKz2RRPR89IHcB5VWsqBBR
tR5ILoi/oWvBCwf4BpHvNaDppltWfdKNdV0eK+BiCN9ypKgQA1LG4EQScPiK+2gmb6dmskKmgfvN
qqUd8qZEtAkXix6y+V6i5ZWFlBHC/xukwbuBu+QQNur/MmfjW4ytIfVxJf46mdcwiN4gHlMGWUv6
zQof4/cNJFcPuCxFwO9NPi/U78uRaOZUj6V1Irtn3jlGJilbuVO3XTRwC7wDQlquw1WUMVVAfbPI
31j7GYKzzIgFzKrbH/kvMZxYZLLQ49+MhKVcAHCb+8UcSDXbwCY8hpM8ObuKSupZmJ6d2PXcr3Tv
2pm4w8qJVN8TRRaubKN2Zh5Q3pofHNrubBSwvsVjlqmqIL4UADTf8Kt2jAdvDe0pJJj2Ur1dZ4ck
myN8esim4LBTSw3SAy4dLYLuCpvK0GeILA/yNg+w+gzPrAjOtMdJZ4Zys4HjFEaFr7Igx9Be+MBZ
l1h1hfJAHIW/bN5TpQhKx3txxFkTadczzIExyEwV4/bqkiJ2nTwE4iGxfwykbKVR2uMMI6AA7jmu
tnuEX6/Y1K6KLWDYfhhCMdd1aM3w4+F73EQzhW4gBq/RfX7hJM4VxSJ7Y6+r3GsD7U5wAu8WbbFy
ZKcJa8vDnit9Q+mgYzXTYKdwCeAhW462tgeJ1mApTS2kOCLTJLlYLmFhgigucK5BONvZGyFUarSG
Ltdud5U0fRUdbduY51k9WvxLF5jc3Sojy4y8KqWpN+k4GDL5EzBnufq49NKnKcDKivRXx3wfBbi+
yMIO0ztE4t8nX/lXyVhZQL5SDFSRHS6YsfeAGBNARH64af1/bXmUQALMiuQY17054ESSRPkOONMK
meOb58y7VKlSsyGSsYjjbEDaJRnxZTnZVbGmTeVMUVDGGai+423Zu7H9FBsshdo2A0oSUaEBTWb2
aeoEJiRfmaG5e4BW3jr5b41ISnh+gAy2M3jF9zjyt2bEMUnrk/CeKFr+jrjG+a+M2keU7cF6d3sK
dLpktNQE6YGtN92eD+pL51Jy6WFN1yUZmhOIaLDtXP7wRy+7+k7259IaQ7XOrEMSblSmHOquqUKB
9pk8fXgrpxV/fVpYNCBP4K7tfeb+XKutYdc3v7hYboNcb80nPDhbAwvXN6fD6kbtEsSmMbXWKMQw
SRR0zt0l718anUPnevuRTvOYJ0C3jfKP2TNwZkoJWNAf/OHc7/rPdc/lLp41Li6vWObzoexKiy3N
qmzkAQzgVEHs9U+34hCSP3UIwnnxpv8ZV7v4WX6e0Mr93A6yNO+q14nrG2cP0vuE5aCSDz35fwEO
0O+tozGABfR4GuT4rJGfHWPaeJ5+dq6/VZ5LCENyYCjdP7xLFcuX5Mwi0O12dFOilaowNdUUJvjI
9QXlrcxPYmu1gPSLgEx7eWv+r7A0Fu1JOvHy835fKPFmFptHOrwtgQo9L/DDuz9JFwqyvR1oqJOB
CYB8PuhFv0mc8FftaSQfUglf7RsLwTUbM0BlE7UJiyXI17lhfCNQrygF/X0PqPSS0kfgHWRWhdJO
gUotCabbsu2FjC/1i9Qa6egb4BnZMnkfP3XPf9CzwVETrv2HmL6i4G67+jifAlYyGqyTR2+ndq6/
YA4LImvEl4Sf0SMEn1Zk/k0wgWNQaawQr0NzmWdnGZtTHuBOR/JG7wkHjImETlSJ98mdmXNb3/Ve
cd9krKZM+3fTGcSbyigqZGDQrcFqUPOG/TQ2Yemdpv21ZnMo1lX2xkxki80yqeOu0sORbSRutFgD
cwQxIf1C5x8k00pzFrLd6U/7dvHGgdx6AvJrSLkCb45n+lWYluUoROkyO8kwwer6CNEDocKKNNBk
Kb2qKThX9Qwo1lfTRy+9n7OzxgIg8s2+8401Bzg5wPJykMXpSGa7tQmmsKFCHnacPJoPsurw2Bqg
k93vJNVFozfKEICytVHctmJhvf+NUETmbw1rjemrTq+Pbt/0FiC0TTOo9CDeUZdj8tCxgFABtft2
jB1MmKsF3e9B/x5dJb1FleGcCtpGkMEz9tlNJm4nN2RNmZFu9Oc1hr5UmJTAZLPwSBXhmqa+bLsO
C2cqyiEtLtsV6U57Yj2t7UqQgCr5HZKGtK+BnOlW4SH482GeHTVSn7SwvAlBjBUBLfZN5XEaZ/Iy
4YNZJ62lkiihHcqtx4bVyuRH+gRwqoz9uQ6+b15XB9KGueGZsAH54KYQr5WRKw5147qON5OEW/nj
cWc/00Dp+AZUhnZrp1k82kTXaH0kcfyA+GYRQ3zsP8odjsa01QZcbX1RPk51WpfKHbkUwDyFCtvC
SRv0xdVmy4BOb/b6KFNsxjdK1E7GvtBV69G/QZk+YPVHdLyGx4Tld9zodxhU8RvklMoRXtjzDB5U
1pU7lrmj/pUPp1Ivu62+NSGEPW9wrgvja594P6Vm5VpmYsee+k5fDpe106aR3p4kjHAoiKRT5zgn
LOWR9FMbh8I2R528+Ehaw+/67fXeEd7txqAHg5qdkGyQU9dDlAqJRb49rOmiw/SUsJfsxLCNRCZ5
YZH9ueH96ft4GWps3J21qzA0jgXwGx6bsvSxpWVQ2dd8Ro89pHoR95dgc7A8st++jaijflaGuOG/
64OYqx95DuO98wIlxAO4wl0Zc2tHwWKMiO6t63StiNcFR3DAbD64vneN+hMHP1rhpPzbCeRZ7v5e
kTCFNuYHxd2EWjPM6UesDIzfZwfgnMP+WONX3t85xqAWxJBiaq6OGCNGyVi40CXhfj6Wt2imaxK2
yjZpzZWczhfPsZq754SmJ8/Lo5dgvM2hijy6EX5RpJhZfpZGCxUsUXthOPG5sk+5Z4dNIubHzivN
mnAflk5Eb8XjbwwmmdbYVC3FtDTvPQ5nPC3Jdwkqm0vXOMrlbzRqM2+Vx2M+5vYL3lgC2CJrP22b
51miq2nXOCkSBuZtRcq21Z19Gu+zcMzQzMxrj540FN0XfEDWPhvbL3rladJPqqdZP/sMQQywgvow
Ymabc7Gf7smmdqKP21LhGPBI4xDlUuzHjj/iBwwtI7iC5lY04ZliVhmDgGlNxt006mlcX5xrGMMY
uNzfBUUtyk0j6gUAG1w92BFYKN5ENPvd+O5iJj/s497z6YLpY15f460Nrnem+cvI4xCE7l1BJVdB
BOR791+N48Pf84VynnQJe9bk83Sd+8mzmhzK5lTm5w3SVIkCtEHy28m5AljganDYlwoNL6y+t/eN
1a04b1gWT/yPPowzF2LtBOUD+K6HzbQLpN+4p8q7CwFEWLyA5JtcwZvlxs5DWeKOrr/1MpC1wv8l
+oOJ89IisquS693H47STmfCCyxZ2FD8My3Sq0fAgvPbUwwYGriE2liiVNTFDzhVpYzn7TTBbbPaT
ZpsR7NpXVQoHVZiW0vp18M9G1liTMt4JcquZjtTdwoyPUzWW+Onodw6KzTY54j/j7Jezqj2744PA
E0erFmTDcn2Y3tOcdzKzgfvSkfEKsAULFssj/HHzgUkV3epp/0h3mw4OHMeh5p/FaB0k6YTAFbtZ
nBxmrq0bVTlmpYZeaGzf7oIvX54BctFBj07ok7FWor9ZJr/gduHhZv/OS5Wn6Gxh5w1h5ipvN0hj
ZkduuzwfF8Cl1upc3y5EEBnsxEuplacv8id0hteLnFVz6VVIO8DCZgwGrOFWKs/Guyq0kwURmNgL
QV6sqIPfkFmo04P6aIAufwE4THkQQVVisE7rGoPbbc5/1vnxA9D5qghaIV5n8b2ZZyvSzOWyNjff
eRXWxkGgQ/CL4PUIyhkjcBiiZCrsTEnidGBTzZohyYMeu5Xx5p5eSP57dvGd1NmVd7blPVRr/8tM
JIDRrkLPS+Bzs55WNihVK/V/uRKatFEzC9AXHyO8+dPWD1sy+qjIM/w1F5aqUh4tn5ZOQmujoE/F
du56GskgXVTLQfKp3PPHG7XVrDQPFr2lUE59a+HOnsDxgh5kYeQoCuxkiQd7ndTu8yQnma6J8Ks+
aS7O9IK/uAq+FDvENN/xmBH+mxOuexWNBY+4y5PJ0LB7+NaDTnrGVXC/BCulvdWdY7VGG8c7/2tc
CF0foA5RAgwANW5XGdQAZ7cnAvLiTx6H5Ty6DUKqBCjJF1gL+hEeym/JXoTEHPXRzeKx0+OMZ6S/
I+vQH3NdT8vFKy9RMG2xwUO3qDds6K3T4PM+l/A5AQYqsBkDO4eMkBKfedADpI7TJdql+fT5LhiB
I4971G6OBZ3OobXrQbibxRydPS8h2FqgMygsZsVGq5nMvpuf/hjQh1Wg7oavYw2jiHIRVcBsK2fr
1pgdvkrbCXA7244yREvHIHPxiuZ010R3f4AQy16dlveAFTWT0FKhLHcjSfdlgGfgb1wqzT6mNur1
gl2sUh873qa3Xoio4QwQOpw18xHtfHuoZl8fznteuZI56r8fWiPSOZtKzz7yGiciVdjiiZe7YWB3
SDvJT2GPW0we3/blV4yZ4sjZoofUodiuYOmQmSl5RprlrLgAtRulrt+n4kreg/qFx3n1A/nv93jI
E5HKb+tTFpKDLSzWZQJxQrg2FVCRGqYFbFdYDFdR3i4KZgQOtq5VqHraAMUw1aLwHeltfs5ltQT6
GGWNnEGo7kQD49x/BSghEb9X5TBW9ouukUf+Ii596XnzLt5+l5tNz48iM9hYErS5bHXx0aSrntq+
LVae/gZP2auhWXKZy0QKU+WWRMLpgXvMYtvsGtjR8uKjKCN1nYI0cHuihgu0b/nsCUoeA9gqr3Kw
Ws5Zb/MxuKpGGKgl9Udg1ZGVgUgItgXBOHXs3o+2rWKH6RS2ljvs5B4s3iQWdvPwqBYeUlKIwNAe
xkr+/KN999e46i3kNS16sdnL77Tlmrye0ZDDoZN00IjLIsRzEfqlEIHMq1XrLKpSL7OAB/frAQq5
5FjVmPVpqIBQpmLA3FlN7Ucr0iTlPg91lIpvHVJRHVnXumQBWWtWbUeueCy+px0DNEEskh48UlDQ
+H0qqC0gzQVqNAu9zm2UMtYqLUaEDwV7BW4XCfUhgAXvycqk2fYcMoAi+WOMiEpBGSYIuPV7pxWF
ZKP9fj415LfCn14ShWktgKO9MJ/3F3QdROD6zONoCP8QT6JkH7+oCJPeaVcOUftJIIBI/fwPiAeG
xKgbJpmIqddcUUzDQidvuLvdloupZuaOXnvC7bU2zIObURMj8MOMbGLkQyFk9o9VHCoKlg50WXK6
z26Z5WkOrEfcxgrdsFRYALDZIXYrrkfKVYDD7t1UkeMTAAUpYEGAWQ1K3QNuO2uijCM4HxkOkOE3
rTSr3FpzbvgrNfEIskBSWC4eS6beSoWMGWQLqNOy1h3+UbKL2cps4+CUrIzYV1zysJv33MkRIQgb
+vF7iU3OAtY1seaDIpy9lCaIjTBHjkPA7/UOrIh0JT06q7MFxu4ksoAnZeDHJB8WLJ2BNP1ovXn/
NklHU1pt3y+806t3K6gNifvUdnOwY0usMqmlzOZJQVSKXJe0nVGkogsxOUGrQcthjI9iAL1wnqip
gd/AzyyRN9tJ0cyWhOZNCFaOFsRPqDu+wMOiaHhQpF2edoEjpwSVLHdoN5qmEZWKMVcK1sphv7Mm
ZCoHHhoYC6usDmsW0LUpMmPNRfF1Szk8OPDMZ9AKtkTIr60naUdGtYLEIk0FiXmykCUZpqL8pG7g
K/7FEwXgrVdt9IwNe0TEgwyYIjR11TwA0kBrXyERRvzsfn196IY4XffA/bQhcCgPfAeKk3MGVgcV
2AFVtspm6bAEkmG4vVFph30tIr0AAwTitJbFeSH95Qxlss/I/OUg8MnITfIZGfyMaoBdwC3Da3nw
5FbLRiQwLun6jaSY+gP3Vm14dh90Dy2r+TG3SkfuRUCmdHYqkERuAq3A/4Fo6LjT91Lc1fqInUSS
SKt5VfrCf+TRYulU+4d0owYvv+W8Y3On/H0PVIDDw5YEs/My2pcHt61v1k+hpOrXJiBhTx0O8FiA
zbm/vIqR481ZrH0HgOHGUfho6DOYkHrfbARCaHN6X14+d++kl4sugecsTnkt+xo5alOAcsJw0P9i
SYGbzjul7tLllOJYq1G9ybihnuA45IBYAM6Ix5P9NRiPl7HcJFNeD1ljo8r/iUUY1vKVyfW5LCWA
T+yw4gbXewjebcPWoLBWmxAm5GejbYCelSS2gkKVf52EM6DXXe/18DG821vtxGzLb8goKRYsUebO
TCBb7Dv8cHvF8zrnoW3pdxYVBtAn089jJ71bGMNyBHc2thgwd/Q5FF12Ls4JWtre2rB246ZJ+o4W
XHDNvAjMBFpbmS3lbmF+tmFHDpARImLrU2HqfcwrDVUO52SuZ32OkGQyIZDaKGwlQgE9fB8WyOQ2
XFIr3lXCQLMBM2xTI/5gpECuTDd3mJ4m9fvsqB1nF4hpXeNZwjoM7VhiWdYYj+Y//40JIv1dFX2J
BOxRDdLal5UR+BIot3RDyhqBJAOUSYYY2O30lONP4azCWyQL9tzMS1PLVCcR5korTYkXaqtq7Ifs
Aid6FfY/m12IZ7UWECMzgZKDcfWGAba/CAIe1BBCV8XAbm7qMTMThjGKUa5a0ICnTSZhaWtYptOJ
O7eqLG1T3mCnvvpMLNaigfdDRYqpdzjlnBnXKJg4uVD4nMD1PEcL/gGxPpKRs5XKkgY99He0YRZP
l8slrOD5wykKsPX+gk3Q5dSY/cNnbjL35Thhl2SZOwv7c8k6RJBGwF2lqpckysHWotTO7rqDJm/U
35ULBqIVkayNLuz/iB8NXuKvOnrAgE6bqFKaaxdTti/vflF4pq31aYHvIYGZBm5nnM9VRuPL9RWk
kiljR6n005gXd4IhKTg1/16nsr1rvpL6GYd0P7WZlbO6w57TUSaonYy+EItixS6xnii4/0IdRifm
HFGHblqbJ3XdTqdbUHHwlWgX6+cm9FXNrhHBMWESq7PIzkDVIaMZcUB7FaYlfY4x4W55GrMjK6+4
5jcWMdq6gzMksoJCqQ28nBPUnZRqiDgyEBhjrYtsyG14duKqalCeNY3LaOHLWEmn0rh9J1Lg9jSD
n6n5WktJdxQjbw70f6EPq/sXmi5wDvumBKPpy6csj8XtrivOAbo2Ep+77ZVT2JZIHFsrSHIxRura
rGsVYx+LhCkLPL36fNrSlo/Ya+lqL7OI73NNFP8fYTUzLNnLZ7961CfjLoXZoZGe7Qgpfx4HqjJm
qYmoAobPOgsihUexbg1OReCukMyutFCRm/5CG4gkciHr70n9u1/4i+zkuR85fTeRpSc7qKMMyCeB
5VA7qf3pPQ9UV2RX2ig956zvmuIGYjStnQpi/QvDmS//PXyzHpfXV9kEgwmyOoUFhryYGcKY/zF4
0cKL37/oJPK7S12wH92XbeBo4FZC/LofliN9YdElYearqteqSnhkgIVx0BsgTT5GWZAqWO7kcouc
rIJgjAosX+E5/sR23BktDpP3HIXb1iI4hbLSK6XZfLMAw51KrAs+uXPUnDXVdJ9se3uyUpJJk120
5oied158L0n/33kCqIGWMCDqyqx/jKI6DrLDKVrP1rNon2zX62KDvgktwlstfqzJa8BajP7eZaeP
VWfs/YQeT8xF39NVFo5uLsnY4R0yn4BaAjfmXLXkyAD+TmuBfkOBziNrH/1DTDB6kasmZavbUBhX
EP9E2/AQ1/Z1L98Pb1xH2N9Tm909/BhqVycabCZ4kKKGYqXXVxCndW1mA2JxH5MRObtLzvj6Agd0
McUPUKWcrKSMRR3Qql+Y4+ZeiRb+i/Qxd/8h9mjrvmR/MHlQS2Y+Amhv81py5cQ2D2peCjXcRE3W
HNNz01W2iLtZfD3kUUEER7XUG3m/ZP82477kBU8jo0cGG4fLZXMCa+457u7MjeJlisNesscR+ErF
pfpDGjJLl7M1N8bMcuuipPz2M6OB7nLSMAZ6P5tNdiAHAaod8xr8K1AfjDJ9mtUfx4+/SMTem7v4
J4JF9Sd2qQfvHGU8am/8OUldR1/7DjYTlbTl/WyLP+SISk8PHpQaezyPTauX4ihUfvzJR+EFTpZa
pQbj4LbwZQCU7j5H0iLW7d7R5Ib6Tjk3ieeLKZ9WTccEQ1V41seZuS07mSS42sADQs2iuiPzYgxr
UOGoexwMY53939rZdhCsH1IYXVJv4fD74hzscYq6KPWtk58eWrRcyqtyanE02PxMYJvHkjpUNvFT
NzeRRvfhMiaq7C4DOgDLoviYE0RTAaQNoxq9UbBl2jjTb2CHNGNZCUG0nnLf74QAc+f20I0uSp47
kEpWbuJWsYZwFjCz81PInRYRn47U1jxAaKHtFzCLVmco4GoDWZsmtVxO5AJ9zss0gla5jy/GKHEH
ozbdvo0XGWDImViaGgWoUoxC+gOpHLPp2958cXNzfA7qs0sHng9WDPS9SZ8sMnlhXCzpJdTmP2Ba
TwUscqJlSUG27FYHABh2f13+BReHwTmUeQSqeDxdvXSwS6rD5IvgSLG3SPFI/cvrgDt70wPVOjuB
qefXMRCIhPH8uyqN+/5nMzvQ0Cal31h8dRza6XgNwukLPq0idhNJYZCvbLDvCngWK2lzJ7LquwXU
VHANAJDVY4m8aUqIItoB8QxYOyT9rWf1eZ6DWLKFkl1iG6x4ZJNJVhg3PXgzQwVfo4tJtW0jjGQD
tzYtHHXnAwJpKueA44JpL/zmfJSR+ooFLQcF92twYy3sqCpWDBadG2jxkwDSmPcxXv/kU+SiZLnc
trek9mHcBVIjZkF03wzyY3rnoaKYXWniS1YKqjm3b2x+nuRhxwVFtr3KVlUSWlz7N5VVqfp2utva
Jj8/1BsCqblup7263nFHpm7h/ZrZn1/JjxU1rPj7GuNYhOb0PB+osnN0eg6o2M1+6Tq25syu0ZIY
5DxK4nqtG64Nfpr6mvrPWHSwDB8jfIavGzmWG1FHRVck0o6MWgkrx6khGR6YEmi11wolPt2a84Q3
k+MAAJzjYyyp6kwQBQ4yFPplSctPkwImzGU5GYMPuX0GD06T9pap6G5zdQ4y3aGS0fgsbNWYRDD5
aHf1UgoMAF8X5lTS8+EP4Dus1ZNFJs9FPXK7XEYvmIJAbPLa8z4ISt7cJypW/8llnN+tPZVOPNSt
cuTn6BiJJi+8AEdIVda8fw0Mz+P79WtBzGZL1kASmnbm4cl4Dsm40dixsjZ8mVHQxd2oIGFl2sTp
FAxbEWFTEdDBxUS90Gj7WMMCANbb+hvEC/fBYqa09d/UhvHYmWG5VfXbjxEDb8ToIZ7QTwBE3Nse
XQ3wGuZGvAlJpygVvdeD0DMchK1kPjrcURbRGs8bwECfbzsRhuKwmneBQ6T71DQUa107JECMU/eE
tEGyeqsEYnC/I3+L5keQNp3d1MB9J0/+oOkPwyp7Dfkii0o3pPcIgUr173YsBTYxA0H+0/yuHCQa
YijD2mUCEEtiDU017KPGczjHzyrv8/Gu82wldlqmr0EYOX7VAncvnTNlsm5xHhtJeu/XXhVW+TkJ
bhzVKi2OBYgTp08vuWikStPdynfHDQmssR+O0SRdOsj9BZxOLA54duJdCeG2N2mhdGQSlzjq5iMY
8UkRzEAIsj1Wew1WFHh24f4O9XzoUOgMWqsSR92aMvbH2PdWKX9KI88Sn4sotnBESMCaKa4WlMcb
5p/P1n8I9b67jqCURIqji79B5GiZ9iGBaOLD7+2M5+DRzs1aJ76FQ1a8DWsgzWPxqxx33OFf//+M
mYO0N+y24rgr3yz+DZ1ZWNDNcfCKANEGfytuDoPI2caMULPzj4PXf6F8qdUnhPQXNjNIInoJtZ9o
p7X445c1M6lZxkry8T2abvMfqnabZlnFMxeg6Z0lEqEV8OCeMp1my0h2lJtSWHRnRTuans0pUpHI
mhdCekumjO3knmHo3WsHWVxeOfVhcZ9mUFMp7t8/F/9+j6XtNJakys+WWjCZ2TxYECFim3tpi6fo
pV+Rjp+WRobnKZEjWZHgAwGtbO/Um6H5GS3tkNuKmhYcigv7ain1wFnlHr6awU4VzrJFPqzK1M75
AgNMB+I04zfMV8hp+w+4tAW4YMmZbA4E9t8Qr0FIixKKP3Kpa9MFzDg3CM2FpIW3ZkmyLiEcYxKv
vxUsFi5XEgUif2xllC4KX9AJ3pKXgwI1cxNguI+LHbaYGn/EUUNQgf44ICO9FF0NWMlh2L2k7q01
CKnieJCIIDdmAhJs6/iGXkgx6xJFXZmk6/msL/uOxCFRXwLfpg+sOz+ol/7Qbd3BKPhBE0Ggh8Dx
4wzgzW/b0aLPhxSts7u1CQOcHoc4TIB7XcMBOXX9QMeTs7qX/EWJDK5u8+KP6ygHURPqyLqZ5w3f
Ut1V1wBo0Pj+KkcEb/OX0vYn7DqQGrzt0kQ+Wz6nVQk1C/Jb/nYNTss6Y1Mon0b94RT4W4K790KQ
Q4Hu0F8zK484R7bXl95+ar2N6RuPd486aFGvyu+Q1YmN4Jk8btJ+dVyUcSDPt7VyAF0YkXYHymq6
GTO8veIM6U46d7KwMMDqi8TEDJtDpROqdWmCQu6yVLLIx1a95DUX41c72VUezyHIkR2eLSqepM6l
ekUArUT4kZ8yMugKW8MkueH0uIfkakQWV0+fvcZxkJ2O/t7T6zzMiRpKWyKJGdNKNLTWaKH+mSUD
QGphsowsyxuOLZmnHmdoyXgGr8Tl5MNTUsWvZlqRtKbnn6d4nE5ypX2P+QCepF/+hcTisW7Ew3Gt
+RIECq/bs4YQ4gUtxPjBnQHXYTOPJ4E5SVVAZbBKPZHriUuBDv9Rudz0HxfnFQ8Kun1oK0ksciyt
0dSJaMxIoN7g08Ll8PH6WBSSWjK26o3lySWCDab+lHb9Zjn3D2yHJHdGVxJRtmRHNVMGO+D1Gtft
uBQ4VmM7ubCuiIbjiD68wx0ZZfH1YIp3VOZvhfMn0sdlTMBVgBRreNFhJxQqPuVIHJG2lpZRBNKp
Ispl4jpimWdkEqJ7mmbKY4izZEioW6xnkgL9fF+eAoGV2Rx/GN7EFAr4DiXaxv7+mbiJ8Ycmi/a8
iYQt+rkcNMapesWl0pEUDnEqvp/ASL1hVhfj6gVsgKcnPLOUSkvXXYoE9d0VQJVa/IRKoA4BXC17
3JxfPCY75fYbnBNDDwXAyxPzTS7lGRF+pDdNyk1lXjml7JJiKa988jbWdjq4Vbb5tsZn9enzs7cp
sgKWTJvaYhYd2NEEIedjQvEyh4vlOjpCq8e4lc5rXjmQ9P8boibYF0Lqnv+oOJGFOJPPTiZVy1WL
VRbfmNfnfR748coRTE3W8pePTKUC84nMsLm7mMXeGnNH7KGi4LnOQ+VZMIcKczBVaNeucx98/+Nl
LRcKcWL0svqYSEeTJAyr7P9C03kLUtQK+EsoI8VFXYQYP7wFDYn3j5BvPuMLgLjTy1SGwx6HfKdA
MA8RuqPSA3eMhWhAdqTufHzLEJ9KHm1cAMYZgjYvtELuug7T6yhkEOhxs/JVlX59RU4Fp+43QyeJ
q69xgLuYCrNI7gvjcRFibYZB/XgIMx/F4SBH6xYj+20O/DytbGyISe6HWzxaBE1305zVKoBBDYfM
P4OKC1YTjvoBln+K1LVGYs1MBLkjQb8+LxulJEb+lD1t7EGhbw2LOq3u1A/OogjagwsYOlwo2J76
TR2vweqnJhb6/fx9Ep3UuBz2MClmYmLGXsDCMQOCGqFHHmtjhHD3+IA7NeC8qbVyl6HshvosF6iO
6CRPJbf+tbB5YjtmvxQ61iTSIDoAiAKbHol7xsA1f5xs1ScLLrLqpL9VO/m9x0CFZHZRupcWHNqQ
P8YY2nnJnv1nc7qR97Uae8ZwKyG0UL/Uz0kxMDV3Ui3Iq3m1BXvF+msF4xjN9arI6jd+fK3oi7nk
ElPZ9RgdJQGx71AY7anWfjwWwIC1OvVjC55tJCEM8VQCUpqyXBaNOOuQZHZzYL+nBbSgLolvtyZt
TXK+LwKudAVwQd8sT0nvzeGppUx8YZR0FqfXqShCKVb93kW2+0yt03ya/fqJ0Aio4z10nZUDOBV6
b8EImJLoaoxjj4iRHXZ2+teQTNYiqGlJJOB8UlY1JaVF/junreuaznx4Pl7YHDRIj0wzshdv1awA
XWU9sQHAwBNf6IqNI7P+UZI6JF79Y+hNTzgm5DPcIwNjrkPu8VIqWhqjGUD5nSIbuv4JOeo5aeVw
6qQu6LyuuikqQMxtyb1WufNNlH8du422WntDtmpEelvIBOn7cgrsCi+m/XkYOrmfXjro5RAF+FOJ
OVl8xiF05iYHXo51GluIj3Vmoti2W1FVFwAm5Y+nIyYJXXq9QRT96uHz7QgQpN3RnkdCOkAxW2bM
FvRKMnqQ7O99EoMDKDmtinSVFYKVIhlI5eFWg76T0AuoaCyKeh6JRgvPcYcWPLfaBCEjUaI/UIUE
9ttD8mrnfyo+5mg/17zct0fobJ9XQ+fFsJ+HSaHn76cOliAPV51j8yT9vZ71tzs0g3ly+bc4hdqo
5NlKNIA4LbLokSz++gadfCU7VKI9qhoJZIYDhzxd3VvGAKp8RX4q69Ersn/NXq9nUqumDbzKiBxv
4uZp6NNU4GecpsPA8P1EIpIV47Jm+pEkqeLirAjmis+BhbRocIFecqEkpgCzO6uA+QDZjM6VR5vy
Pc3/xXs22jwPK+X99+qnLaS+VeIhBoxgE/i/Z4VHOHdjBYskxQFB9A5hf8uHrs+VFaVpjfrpV9l2
5FKatTsFZAI0WdkFbjC9txiL6o58QLwbd0JahqZt+kPBTRcaU+C0Yr41v9jZ8e1RPHfCUmf7qvD8
xdhEqYVQB7jC8YMnR6aV+8pbraKWTfpBkHimlXrs3dlC4Q6LXdaFgLjS8b5FLU+62aXq1eEiH13k
2nN3hzj9yP5KT9yu+pWgjnaA9JXgSbgcCSX3n10EMjr+3h+QtjCXsNNH9mxCQEJ0vd7IFGA5BjkO
WWwNUSkY/2fWU1pbVzvsmUsPMF4rxwb+MOT+CyLcTqQMMGZgU+xJUjctivXc+qp8CRzKaQKVmoXI
01t+veHVb9ul8AFcgr2stmBKhTtIj8ggn2ThbqOVuXo4/jDMU9gQtDeO9JcHrqHr4OqYQdQzYmQV
O60ubSCfAkeofYaEDlOkrtZkYSmNc+yp5XvPwg/hNnSW5E+RHS2GVWcY/M4IlHjrx9ViQBVQ+1/N
Q9ikgKt3sk7mlxjwULT9+Dsk6kgHAVevq5yyJDmQkIBdbKM82FiUM+RfXh8/U728SJRgB55XdwJ7
t5zvEG33hsPEU/NgxMAVw397vp6GRVwteFxkBdDOtXf1q3W7XylEerYhwcpdCoRh6PyMkTxlwyiU
ld9iRq5s8G1wDicSSePDMSzmJz6tkVLwr5WZK6M9tdCy3YNSRy1+JuCy86Ttd58hTlZ+w6HJgWis
kCPHnszYlkyPj4LW+35zLY4X/4dt66HtjxuS3XBAo3VRWUO3AkF4g1jfFDheV0LksOnjqosRXgek
9DvmooPVQdcXqIaxMa9zPO2XKEmVt7/4xVRmFWW3bdkvTt096p+wfiO5azvisE4q4lCub5X7fiWL
ewOPDD7iw9t7ZUBgrvsUbZ/YpwS7CJECO9HeeudMTr9gYkuXocaicgJEY2L0Tf0u+6ojzy6u+K9H
GPrPShyXntzfiU/9OIhW/3rrKvcNShf8h2oQkdy5H7HmdzCNV7XUte56o7QSHQoXPHrYa7R079nN
naif2YL40GCfqgi5n1hk7O5TCEGU/WcBlgk4y/juNi8M7oNlalyyNI7mCGQEkJRA4nyGAr0HFdae
VAjXMsmmn1ILhglZrqvMiMRJtsYlhmQ/Z6AE1pyO7ljzmRJui+atx2iyTnUEVqIHa8lw7/yhENqb
tQr6IzVSmCyEmN0/zNx6t+deGkGqDG2uPRJ9/6isYiA3+6/q1TeuI6p4c7KLtzX6nyg5rFuC7j1k
0y91rSP6KMGhSokzW69fzSIF3STmCzFtRdS8e352lql1PlpYxv/6Xi9Bit+1752IynOuavYphmxD
m/MIjHYp81Z8oKW3Y35l1y+PJlp4yIKN4LbgkS/7bcRMChOURRBosZ8Ti/6SxzqlHk5i+givxUCe
FsyEAU75bfIlUabim6M4JpeWBNzpT42D+0+53ADOGUvz5CikRzk9RLR32tf2RN/vL600qBbyQhhK
SuiBzw/EwcOIe17AA85cfpJ0Afgrx0c7kdbKvYsEpEcrrAS+6DQG43oTH8drlXDUgc5SeNOmHHAJ
bTOg3ApUYF1e+bnyj8/jOhxESRkhRSuRT/Xy50oyVwL8+GqZN6oOH2HVsJBs+Vu6eDD7vtidT3A0
uM3o2ugl7bTiHBWLNlAS30IUPacwRBw5qO2SZrCPIYs8fMIQ6AUdNeXUUgL+a051cO+47HGH9ASs
4uVQgJBWzGy2D0UhF7LyrcZfhSVRD2skE00t7VPNIgzuAhwc5vVwVZPgZs5dVKxrE0F/pEKVWORH
geQrPXhECuRwjRscwhx9mxBgGtOnxgRuoGPY/Ai9GSCsNDagatmsORxrh4T6uFuZ0xep8FQjNK5t
q4leTNJbNnAgYO9YB5DK4uQCJmcdTtzvm40T8yB2VcjZSrRD29xuA0zqlOCpydpRataQAGd4E5fV
tunaubY/bCRaSyTasyd//1MEHFwIHNkgfqW988d3pXd3lPaMQvFMb9/w8buYLplDJNNLBXP1n4Bu
ugY0YEzgyDCntSmFcODZ0k7jYDmB418FxvefhRYUlSJBuuccVvL01+JQNH9q1OApnlE3Mlp63gGq
1v/ug+HBudHs0ExequV/l4GZxjfeSz8w1/iIJqJjCZyZc/oxH4cfrzIObkyx3PBkXETHDQNlA99l
+xpyfGu6IN0iIpo0cdqHblZnW5JuddZE4vr82grtbuO+006Z9Rh/hcZgQUch1Xr3RzoFhwNz6uJk
lpOR8ZDe5ylAO/jF96giUTRbUZiDRBnz1L+IqIgr8t8H5n+1KLd2Miv7TCmst7RsUY9LXsOXgv1E
kno2dmzQbQCY5SETyLh9lfZdJPJTghyDXoIuU+uKkqnTkIf4Q8t9EC7okCBkPccga45Dw0+VOEMk
AZvkCsXluHwz8KitYI1GfXEKDXkcZZl9Kp0cwUHubso+hcAqS+sy6v5hHrZeYFAXKc1VYgHNwqKn
rPwjzNyJzrYmIlRQsqU+hnUTz489l+9aSA+spcGvVvZJugj34b3qQ914HVdLnOANnwalIoSL/8Cr
xX0aL4J0aO14cWLu8Ml9hMDmOKtAqVypqWR+IH2UQkIspJVGZbYa4bh1LsfMR57Gbkas82f8yd9C
T6TNZPUgVEPzbXdwWemK78MyWEzafh6picaIa+nPjNUM8C4Lh3NFS3gp9PGGMDMPjzk2lnlU4nj3
bi5jRJq29jx+bx8V46aM01WQgilWFesDpdlgKT06JRa4QEi/KrQV4qwJAxjb9Db2p7UPklvD9JZf
4CIS1qRm30yq+FjFOmmpK4Py53UNtj86k61GaatKfYAh8BN+DChbjxhkpdLpoL27VfoFlwZ5ttso
4qFEvL5dQ8EEQmtS4DQjdWhWI7sWLB+26SeABAJrQNUEnoui/NQlcGZfbZWpw+LQPOvva6+PlZ2P
Y2oFG6WzI+XOnaBliRLQYwum+4K7Cz/V2F8Ih5inxz8O2alEre9EV1kvJaPb5zzc3JejaXOZ0KyU
vtB9Mwt1267PBztlbaDM7sQYOHl5y9z5f2iH5Hj/JIhIR7Qk9vdoek1/sRh5z1+G58CkXReasGSm
TP2qQo6xieIL2vSulzaJxVrrHviAaitUAiw0AOTa4Oa65j47iMuno4B7+d55tayxfQddvFWBAk2d
eAfl++hIeYmjroJAUyL4HDAwgKv6uQTe2u+lLxpvMVz0m14vwRwF5rifEmYX9fFNGKd/e8X/tXlP
bawQryMjTZgEsSeQk5JrY2/B/Q6wbM4i+aia4aqveHrmsxfJX7p4OOGf0neg5vaEbl1Y5AMCpyBX
KM/HO1xRgFuM41+/Mkg2Q8iqkMuTqhBdjmvM7wG7i3fvaUU2w4+36OF5f2oOab4Fl5zWjYig9VAO
kBN6il0poKYqFzxAB2UdQDRRgLWlm9KgutawgFNXxh/ZCtKHyLBeYBtEPMSSn/qfokTgSRT4CmTE
pjMyImlQkIgt3NJWlr4MstCLAIL1DvUPfLu/X931Cr652+fDrUVvTjTvL+1a9pdrq78LROV5sYpP
+UqN34gkaNbph+op595ZT4ArWw4Z+qiZ5bhAVUs1HvAfO8WoRxmZUaCw4cNgmQ6CAYMGkGZHvuPX
qPdL+E0Xoczutn8vSQudv+sYiqLHSpbuGbDLMscYgVUyLK2i5nzGE7N08vlL6Op1oVGcykJdYLm3
Zg/pVo7loyejZu/+ZH4xWrmBB6LmLii3pxr2sPqbBQea1+i3i46X96WG3ehL9KAeB2SjQwL4iqX3
ppjJvNvTnlyM0+LrIcTMO/YQfP45vtHr89ZndcTIg9shi+8KK0pyWuVdzQicBA+Dl9pmS419ZtPx
jKaktloD8f1GrHH80chtqtuz0ZYO0gv5io75UVAjPbINFuuACi48GYgqPXj6aSC6RrgKc8ZENumD
JoYpnwBOb67HWPfcfSb3goQiVgCCPcHoCjVcT2YlVeW8CLaSK3QMMXT6+Q5KLDHG8ETWfWChbal3
C+7B9GTY442/kM0fdG+Xna2p2vqTK84nr4rwde4dhQo+y+wQDSyTRYeCCisgwVLsV9NVhIdQjDOl
QYmeOFrA5y8tlFoJnQloScFrza/DpXP2JeMI7jSJhnPTwKX71JyQRuFgS08xhz7gycRxtK06XzjI
2qfa/Nw+0njqcIpS5M5p+1YWYEhkh/XhHmOVD/xbN7iUNTjgCEId/k3dzh/mJ8NZFY9Sav2O+Gp2
EXgKZjK2B1pFAlgzCFk8EdFxcVzQPLs/CCguj1TSf9pzU0cA36fvprAmQHQSrVNnxgqM3tHgCvSv
ufmVrOYfPDLvw9bsqq7xOZQf3PHGd7Is02Q6QRxFiKCo+QsExJsc1eiTQXp376z3+NTHxThsPzGL
SE2Jw9BzNgbqLOu2ZZsXRaaQGjL/S70g/x6Lt3QmkfcV77Sbc/Wv2TgKcoT0wDLzJOCKwJLh/1R7
Z6QHkP91neNrDIK5nqUO3sOIq8frMObbfKThMFPBuogp2l2NFl1kYjsm2bV68ZPSQZSLa0YVKqlu
xNbOc1Cfs75nDyAVPKxn0muqhCF3P2NgHQnhtcdp9ssUyoSClhEvFB/Uz95HRxihN2ZcAVH8etIy
tk22c9XykoVYkoSHqag8yMDYv4k2wDgmUVdfULV6zggHYfL3/YMA1nom9uzico82AisGUo1C2dhF
Q67RnfE7OPCDcfLtluAD5NLMZkqtcIjFXPWyAvceO/x35G9b4jX4gSTVxrob+tHRxRa9GvHpQJkM
EjL8GY0WYhNTXJJwQTsGce6yD/KSjIQ63CZ6Ev5oR/MD7v/7CPWGB8MbUMGTrajolK6xS8uzD7y1
KbaIKAB+Aki0PDv+aRZOnv9ZwDfLLq+828lNBW7vkF1yH4Nt05+DS2hcFhayeZeog2fDx3ccVzMr
63xYOrJLnz5uwGzvKijgulzc/VPJca/2bBS9Uhws0vu7tJs8C3/z7Y0O0z1S7cU9NnfYJkw/77Qy
g0f6qUGBIcbbY7gZYexa1UJ4G+Hd9T2l2fY+lgBqEvKTzJXTxzRMYm4l/x2y9gJO5tOBsgcruNfU
6LOkvSlIE02M/FCkUTgbmiLe/2flyf9ziXhom6ZroUvrz1g6XPrIR2syyhepu8Wqmq/v854Pzx5E
6ij0SqGriT5CTNk5LOa2RrL2UOwxhhuVp8l/balO+D3Zn3ZZOU3CfYY8aLTLav2jMTWP8w0lej3i
LpFWlFzjIVYX0vTjpA3yiyN1IR1Mqd83zQdaME6aaMll0X+AoQVB7tY8UUdgQFNsBaylR8mqbszw
Zg0AEBV8xty+kckph1Cne3vxvVga2sEHvM+x7/tQ/GPBNMlq/a/6EEx8vY/15j6mWI4cGoZIRyZ3
ejWQ802BBa6I2tas25+ITvrFn+hMsN4i8DUfN5F0VHzJxyNkqqV0Ey8MbUR36Yd94bz46ehzTH+0
9w3twBnmnSIktbwXH1QHaxIqlQy6o1jPt4luhXr2xddNxOYnnjROjrv0KegRZPyHSmrlZbySKcgq
p8Oz7BwS/nnzH2uVe0oVgHBrwQJ/AoHYop6qJOw2vD5IupEELu2VMYdNVVQC7DGp6khd63H2LW0j
auDfQSticM2hF8ZAXkaB3UzM8K++c5/4RXybKK0UdWwR6ux8J9FJMkFKr43Dx2X+7y0chS1nsEE+
UgvWT8w7/uJjd5ADnps2ne6lFmciX89uAiqybruJygQ6LnTFtVpYaONDK6yZl7PrCyByeX4t0Dfx
CC/JCfr0Q3faJEvxMiRxzpI1/+vgsVh2XKUMNX/m/a5u0HyrQrwk3iFfnuiz2vySfcq8jGTBvCiO
RfVIwgdJw4JEJSJDWbqenJT33Vh4qbCdOduXy6U9AwURvi9dYJR4UgUVVnLxcv61FdXLXkH/FP16
fn2IMsh7pJ17xR0lwN2yXsL+ilfe2fLJRNATGvJFoFCPKdJ9fSOZ+VGCPc8o3UP1DmV7oo3yFebs
OXlVkxlsOiUE8cyUT67sYfY7GDliHiSvSnu9vS5q6AEHPrIpnlQYezlWiwB0tarA9RyqUKVlXils
kYJtpxMtSpZ63CDnxdVwFWai8nWILywyaMbOe/w+hKEKGR2zeq2RZ4Ieq805GoiuqanW9LUV80gf
amw+Xe1nZH1jNdq2YyhW6AHXTZN6W9doJQM05zMtwTSRMwwPTBE9xmK0PQh8Djtg9t8sc8AQtzCr
d+hYNUuGd+Vzf5TkIpWMq7+YnKbhSaI+/oKRAREHdvZup8Ab4MKyUsFj17HYPVlcfP9tbmhfmHkN
HtJVq+QQspFGXYf851NQsbDO4z/TQpbk3P8Ki482PBTDbg1UawasUV7samQrqEtgywzwzRWpfswy
DK6NweXbVA3jN6Q1KugLWeBUrT4/e5/h6QCzFn70w0jJIa3ogpuBQeZmAAIcJQHhe9TZkmauqLvG
C7UJqL5zVIRtW/B4ZSIOkfIR9FoASaY1wbBF2rlvtV1owyaON1rWEC3+Japkxes5kIxjCVxLBEHD
MApTjD6gHWHSAIo1i8LVke5OnMGxBig0rTx23Cwu8TzlUeeluSarG8exqhI4fz3FS2kg77A8axoZ
vj9OhHtqYXNc8Uhb8wrvhZBYN9ay4c4zFduPm66qZTrCEOa2B8g+fVW+WohOIMMn9YO/Fk+Eb+ni
QzKE8QNaMOV4tomTetDEXrBoAl+C8xaDfM+EbactoAfdzjS/wPdTE0CCIFYx8lPaYVe24UVxvifv
6MX/IwdFtA/MwfvOX95II8EnEubwaYYDsTP180dqi/L7pdYXziXsBXDJ/Thz1vrb/3x4tZU+W4Tu
LRpOeCZHU98h0xXXGra+I3IKPboCOfH/pqus5KcsbzEfr4qxMSpztXQ6VYVxkP/OpdrGvOklQa4x
PFTq4l52CmXWMKDnW5FBwqFMfi5XPTRu4vwZmBN6Xco51HgTO0phfLqwaQvASy/Utzv4Rxyokngo
dWnuuN8s6ZgzTYAoNbFQ7LdnhfxBY2U0WO3wHFgnO/6w8MhhOY9kL0N60nspDSf1eqbxY4YQkIxE
a5dgcE/Z+BEa084qubZ6K6v+FiaVy89vw3BMiIbwu/ccHx0QLRjdpCSEB5mpSgK3/l0UyomGdeDM
iRW8hmwFSBLvgJNq76ubxJOqZteJ8HuQcMvd4020pIdsLTKBI2snTwZvED2cE7BsLPuMNxwYiXrr
8FJYnP9sGO0by0XcX4yb/S3b8rPBZT1B9iDdUSQz5RsPOHLKKYsCs1TpBOMo051EbRL14zRsYpUv
qm/dHXtfZGzlurLoQQTcY4KWWDKGtV8O+K1GyvFwka1JDMvWmWfeoT6Bgddg8F1zigPwT53/527F
NOGm3TecGhtQkXdwfEowx2PI4XUNXSXngVM0wQ4mRv0M0ResVa5nmjuJIptqURoDxgMXD6q5KjzJ
NrxNqJzhZtE1Hp3nLQOZ/8kFsqzPiRBN2vko9BpFgSCzp+6IeYYtukKnAg53pO3tHUm+kEO6/aD4
LQZqSRENj1Z4xgwCvixW2D6DIplK8fO56H3vSw875yVC07pAtmG+l5j9juczqR3dY3CxvLOBwGz1
BGNzIhpOGD0zAy9LwqD7TnSvnS5oruxLeLTel5NzmjHKXzTWhOeni6poZ+Mu/ySALev5blGpnG41
e1RAl+XmlJGLVcHN8vEMGdTdxEvfyv8FeSdQByjZ3O9S6tZ/YIfg6zzmaqhzNfL97KItPr6BZA4h
JdX5RKfC+koFLePyASJfqRjFTM4uMwfzdN79xaR/mrPcqOSsmXqbgadt7LmNgO3AhOsFlW/r58nz
SdO9FljGQLnH0v47zKnIIjexvWqQLLETMWbreKHlkMqr18BMCEI+ND1VVBzby222j5lK0geapkut
fmqHH+LfZWwT4j3/pY2XJlxHGiAuj8hSdKUgzF7rS7uO2ycBPrz+0ALXw4UW1+NTCxDIkSD0rs10
GeOqkUs+EypIeKuwZ/4kn+LjmkN03S8QATn60hCbuljntwuOJfhO8INd92OJ0kJVuMndSutqFuIH
qsxEvNp2Em5SO4WXYbFKiFOab63IGFfzs5+h3VkAYjZ1GiJ59s1nX0HNZodgo/WMH0JoBBxkwv3w
ZsBrE78/i/DmZFWE7NwduZCrz25kPC32mz4Cwozw1YeeF3I7oBJ6+xMBshd7saots+zACPSjkm0K
rBJs8UaWU2mp+kM1CTc2tMXKPzT+QS/ywZ1skSh02N3Ddq4OVfCzp4cDodCP5cDHrVrA9BZ3icDQ
KU0HpoICJ46hZ1gQDvxsoNoJ9I9sKc+jIFvWVptsRPE/Gqmd7hmB7VjhGW9nvvtcC+buzo1rIjOj
0gsAl0dO3tt0iqe79Ycu9FLRmWn/1EDl5BGPkzFNESH5Dhf+F7dZnCTsdDvza0qJezC58LVu76Gq
G6FfxOhQchpTHgwjRJjIBnoc4sbUMJ+stpEPuDrZ+yJkpw8p2T+EGPP1zF/VhhABbVl+jO3wMh7Q
zh32AihYwEgSq/C1DB045y52b7P/uWiye75cF0d9fdrqu4Si3t0sqbSgEOTANew2XdBicP+SyIAy
w+EatxNt6jb3ojPMnmINHQJ6UkRTZrrRtrDADK45PmbsHzzcee/L13ggiXktWBw28X370ADpnvrH
PcekTJwMDoAnRF0Pf8T1WDjL7U4+KyHq2DyrqkgWrR8WXJfKZC2QZFIg75mg/aZOuV1OVvur8O+U
KIXO1+slPuTkAWUnOutYgb1EEhlFRu04YLVVKVu7FzS4b2WHfiCjfImVvTvvZBjN4Ygheq6a/Mqr
txMMp3nE5AApqzZ/vgzXgY8HV5Hbrf8PKm6Ldl4Mb7CjH/cv/06VS6cOguUw79km809yDbNZxyn4
wfG+1qbvKDgVdJSKonPcM+9hznJpIPRfhTse9E5N1TyZLovE81W4mX/dtwt7pka9msDDq0A9vhbQ
oyB9lIbeGPsYCEyLKKl5/c+B1NmO77ifvThJEKgNj8jyj3Hskob27xN2IRbdnulM9iJSdUqpWqQj
KW2zBO//So+CliS1NZrNn1MryZPxcAj0N9WOwd9HW5CXSMgBzpb3fDU4BfnuaN0QhXK6PA8evY4G
v4eCWFAll491bhfS4TwairyZF05pSyN1GpesX3tnrgGnr/yngJ0UIOKJAGPY5r9JDuUS7zWbjrGX
6Ub8aOsfhM2aW/6CCCCftiwK6JDfh1HN8UUkY0zqti5nYLMZr8zVkbwvpS4Kx0Mq91X2bEEYTvtQ
BLvny93CnCbmxauHG5GQC/sD0oghIFoUwI24a7lWe+m1xQvNwF2kHd2E+7Hj7wTlPx+hIITODXMQ
d0zjW66m+3eiXBc4Pclatiw6fBaHrEklSuPqBJT5JsLVrzoVrmPmPUEEyuJO9cqYrC/+5TvQDi/L
+7/ghs0IwBRpE+ZusfrG7cdJTF0SucN3dNwErivi9ZDwRFLYZ63Vya/bl5V9qbdKTuf+xWwD3ZxH
umWAqxBfdyezstzPZr4E26IZEz7bIpwj5sa/UfHTjJP9XPmqsj/juMF187PruTpD+cquqp/zPT3h
r9KY82EEJcFUt8M7O/Fm16aIPtiRVa70I6C+bN+o7BO2m6E7f+5RV1XOGbVUSBSSYlp3LK5E4nMW
tZR9Q5U0C7H7tOd6HA+mjxGTxuVXmheR+6rqJHmWvjrNhQzn1YVPnbC1uMW+M3YmY0UtQxrY7DRH
6nDJk28oRzl+vyF3Zj+GK4RzHR3p3E5qvyn/W6ZAVPa7qQXCosVWqC/eEZVeK5YtE844+JWczyjH
Dw3ptMzIVxKde2CkCmeNWUJiL5mmMIs50YAb9vLhPdDVPO0AkdHdAtFEiSokGXneX0eakCykc555
/YoqNgTxOylCcE8NvYOksWzUNVaLyncvWRWsiHcDQHmDMo6TpdAbepkuy33V6H2HshMLB0i2SX87
j1iYEJhO3UI6vU+CL7LP84TjH59iHR0eR20aUUvpJn13YUvjTWaIfYqHSQ/Hvf8FV7r6ggFVbw6b
YK+IijCsY+mC6CVkKOzQNkzS7TEUUHznWSYtF2equyaveMVTV3T3FDt9rMOPJf/JciEQjrlUvTny
0vLRdGPLc0Xh99Epr9qpnJpHUXQjSfaIgWWNNfZyIF6if0DUfzyVW9XRmveIclvWwJgj0ddh7Oy2
D536EkxuRnf4/nx7xZ/Q5wMNcoyu7Ht0Ze3hfv9O/0vjIlWloi1xrGHBZzJoinqRQSHaGs6iFJtb
wUpw2BaSl5ObXklllwoMhLNcZecfw9mxkp2XpF5ez/JqN46ASw6/VzT3+FR7d1qFgfkAOZdIDOB5
U/W6dTkTFkNzTN0VrFu6rwvDNrApDcfhK/parIOYlgctw78T2jUJFQ5zXtFPuxZ74oNvC6BVVOOV
JlJl+2ZbDxuA61G2N8mc3ZAZxDywAmjcJlIpEeqPl5iErdXQy1PS+0xpRih7x6G2/8oJYrBx9vZy
3nOChsrp6d45SZxDiu07KK6HDEVmNaujFTRgPNjaFr1CivUeea+sx+fU/44tFi1PR9l7udxSD+XN
HccRA2svfgaRIj4EInB5z+xPAHJ5IsuEQBfuHnbXu/YaUZ8KzLJQbjRX3vuZOLedF+sNLp/uuBS+
7v/O514Pk6XJVHPVQNWiQldyeEB+8fjQsFSzXB3OHyxZfXvDyerK6Q+lwKweVCtWYGcDUZGFZm7H
0CEHT1x1TwYoukOmBgWddY9/fxiN+zVefnVdZwt0UvUXMokxdfMctFM/7M3yMY/Z2c/SIjNzbNzl
3wOhbB53pmYvXbb2T2zG9lyvs57p0w86CRWcqEoLJaCBaaCUsBjL+ZL97azy2mS5/V4LYSvJb8oF
CoXl5VylIwwp2Xs4nhBVoMx4SbqsVPecgQJcKSS0Kr07WhOfStFxZGVq+DroBb+KpSqCnZDn+uIQ
6t+dDbfv3OJGjWw3o1x1cAOKvnn2WR8g0f93hf4A4TZT8maGrJJY7ZVobmsr4IljfHL3SnuceyPf
AuBh3mguOxeKZWOh5QQXLKdbVklTmy44w9j3vd88OWxj7I94UFlrRgeDzjap6+nRkmUy8GDqC/Ax
g8ObzVejKk8J287p/iAmeRsQB7YCDf5pxfwwL6A2R8LBWo2y/NF0KzAEKae/tYpZnDZRVugNYeiW
BGjI3XGag99Jo4XtK+i0uepsp6ptSvkw5P9bqsIFrC7kXjwPOJTGyOR/ptY9/ZW2/mC3+04+OdLu
xJqbQu9Kch2wYoaxAqIEt4Sd8Y6+9nIm8Dv0L3qJAmnyOsDRZuuevYtvmd12mH/8gx3BE56bQo7K
vMtlP74N4YaJSaf4IWgwKyu5SuIenBDkRvwYp1XPk+EaKqvd8uzi589N70gfnFFU4FtM2tLR2dzo
VTV+RfMDRAEW6ruiT+gR61i2qqzeZKNhIuFnDBnkL76c7etKdVbMNODbParvL7FCZfB8mZLnxgYU
CHufQzpHEFYbFZoICSKFNiNZq4stAsBYvVq1zQek345Q7yH6onZlfRrAmpEqLcghlWXdJ0y0Q2ur
fXrEJ8DGeQgODXaLEv89bGEufn3+YSeXa7NrQ73KP7MQcxGcV8C3UntyRQr92atTz6xfGdi4IhRd
uQFSoz8Mucit/mP5yNZEzjOAklLms8MUilvaGf4rkzxTapzEpLVb5QGCSmp6UfnQPS89p1qbT3fN
0noNbKfTXztHWvXwIWbZ/boThn6HRBIei7WS6Q4WgmHMT1Xnns2dL+mOHdRL2e+BSV/cXSb/kjEs
/gGyHGZDrplPDVxL4zhayAsLamXTclYX4hWylpnc54qEyIPVQ2ddYMJYJP+crrVnz0DeHJzDDSjo
WWuDVQvfZiIQmp06TRbZiLIifntnTXstFbH8VV9VMJBlIOD4BbcBaNtTEbBGxYklL9HjxCtf612p
y9jQbjLzRU+y690SBo7+38gq+00tn78uTYxZ/6XBiU/Gf6tPy0F5eHSShr2k6/1NQH140g8s8gd7
o/v+xZLzOtJhdUH2Mw9TVUpctBlJg8Hc6kgWq7u7sOcTqnga4aqrLu3mQVyu62tiTB4xX4sKU5Wf
B4PeeTGFT/p1SC4fEKrJ/SRzW3hr2N8QGjaXX64W69oQMYi+zS/jXIcns/jzU12dDJJjvSLRRKAr
2bK7zmJrvuAvkCFbUSSp39V6j/H6TWTjO9GaZNz70aZhq8AhRUbO4NQq0Vbi+W7Tf73p21xpAkYz
81BdZw6JJzfWKupQjKPQQnlUCiKWDOpONXZMx8ZVsd481i4Nfoe8n/g3stfRfkN8TFXTuqeKENSf
uQb82yUI+tDUrS1FOhvRbyDI7MM2MNRwYWalGlUxUSTjd1MAKTdmTfuzS4W+nbhBGQFvMntUwcmJ
iK/8L+SPb40n0yPZkSUfMYavk3f8GEPzJQfofgbzUqqgrRuchz7Svg606Hg3IC+oBgyNg8w+qjaH
N2N/00YEFH2A9IPA1uqXKagOwOOKpxHyBSjvsPnAQ1j8EyXfMMzQqj1XOYXgQLXCpfocJZheRB62
TgN/LmAbed46xeNTtkRk7g1fCxpmOME4IzyazX7O91ohgyrqURNsbB86IaLiivkL+vETU0K5Fgd3
Nck7A7VsEXDU9hOTghzAzDEXFzEYxhiBQGVuqzGaaYze/ilXrTPUpDxHoBaQu5hnNa9XfDN09Asg
E9rxF9eAzE3CweV15Gkcjo2ILojimqFFZ/AcC5PTmFspC2x5OhXv5XDyhfJ6OkyhZEL64ail1y16
zIUgEo32CLmoyCWNCPnQ9/9PukJj87ponGxxpXW7yarN4vuG4QJhONcw9lKbU9Y8kCsoXTgfYMSl
q4ZxN/qaFiHituYqi6wb40JqKMHgGY7jvJhOjzm5L6NE3cH8oBtS13N328426fyWsR9TNj0SPgpb
Ht/OwYJSpNR/Ie90wf0qTtQhS54hYVE9INW5ahsPdpv+msaD173rI8ea7js2rxp1q31GKZZaDg1X
noiv0FMLt2jVKD3gSvxLG8uqprbOU+o85gi2MFpjaN9ygnr9CVZsPu9S123jVX/GH1RCaQ/Eq1bv
HdVW9FhWkvEDu/LrRCYGpqB73WWU/GZ/YThw7Qtor4hwIsXLL652hGgbWw6jAVx5jYMtQxRzZQB4
ral7ygbdNi0asqiiH1yh64pF7L7FYRIu8z1joVt5hE5zBB5LMgrqD9RuY/z2tQhj9wIeCSC136dg
9tGnf9huRU1MIHchos/5loisv6+Z/pOGl2X98tVkHqyvmX/5q1rIzYj3FCaA4eo5P40h4IxbgWxh
JFBoXmPac0BF6E9X2sIVn0qfZdAyFMBHyzD6/H5P+vnYlKx9y4QwJ6bUcjOdyi2SoS6wgP8vnw69
15MI5Zn1/ZbFZm05xuQu5UY7l4AphW3S6LBIFXnbK0n1baM+r1MrEAz59QBOdZMYxMh0EhEhfiqB
KAtau7+VZbY0W3iWN26Q73ijudoe8e55aO0EVLkYrAJRbhpjuQjyg/3gJDrPnAoQVb+/roxTz5SW
gbOOqoQL3PhBWhM9+2FVJeFSAWMvI5nLoaH8fPws3kw8aJcuMfVucfvOfKdVKW5Fr4B08Nd4EHo3
i6/vzI+HODEenekPVyT+S093wnj9FqqjengxbAZVOMmaDgFt36e0qzKKEGyLo1xxjhPooS1mJeqS
juTXkjGbWkzjnovKM2GAU1uh5e9zXtzPOUAYo5+yVuLLfK1/GLLO1R9iT8wPoFnIRfEaFGoQnDul
Qrnv/+orfLJ0FDRoED4t34pHgcze9F3/faiwdRPbOISSA6p/TiOQVTM5cp7U/Dxshd3cdZ7k71xK
OsTdURQu32InTTZKd9Z34zGhYellUmJn1WBEXM8gdtiAu7bwb8Qottr24GGJoFiVyOKNfEDqqAwi
aLUPr3H4MEkXvI5LSJJH2rHFPHVExfjs9IoWLNrgLXE5hBx1dzUfBvtKmegISfz4mF1pk5PmvxoI
MQix731JZTvfzaOGPaO7HlZsmHra9vd0Sg1lbLT3ZrIvtpGeDd4kS9cSaVENBdPOYklzWIaG57s+
cPCrX7TJr30REY5B5G1BowiTS0XnbxZoZerRn16mTAtYFeZnqe5sN0gQcu1krWhV63vtgrt9UH5M
eLeOqztX64seamQoHdK+F+n/u/PB/WqgRLd5w1FGoiw5vTRL665VZ1kBmNObI9QjnDu2IIh3pRYg
ZBgmY7N5h8AyzlH1EEdICY/sd4p2kpv8Scu3uEbRqf2yWUuPR4fzWWsfva4SVZA3WO7Y2gLgHB7l
h2odtqDn6wYx5Y7ciljJZnyCt8HjJrePKU3nGFstmh+DjnaVcatF4GYcC3r5IFzmHLbrA68y2Kal
szFsWljK3XBP2uvLPcAmNMHpnXhUbn/8sOT89W+aOyYXhPxE5J7PmaC+TEpf+KKcsE0XYYTdv3aD
7niPfTcpqYkO6e58mjcmHcJVtT21Qp7Xz+FF2cXFkgUrvdghwsMaHJ3DBvKT/KlbkNv8QW6P2ax2
IxSwD8/WdIKYxXmvLezAmIkPmFmZGYt7ptnJpz7/oC0AvqGXoMC4Gy0mQjOxJ4EF5RS7V3QLK98i
lkaz3Cf5Wpv4b8M5z02K5/vbBt8T3PnjPZG0IzDTybutpaMy7mGVrRZMpIU6aJmX3xMsHcRniBQk
7X3/J1oGcMLk9M1GwBuFKIIm++Bj9A/iFrpdwQ/wmaU11esew7UkVdQVSszB5Sgqq27EE/RUqq1p
9sqUvq2PhlDXuY/ZFkHi85K4LvIqoCnRGu8fa5JN7TQ2jAK/JfEIXc4gt0Ri09g75kRBiI+tlD7d
dXL3SLIeM/ScIj3nEG7NSdYimt4iNGdmq4sF0KN2rTJGLxR4RKYKWIGoOssqJGYuni6p13AFAGUk
wOVXrVgz5IzgpV84W77TbDs00L4wXIu1egQf6L+yl+0lH+D7+6UWlo1+oV+9Nx3fLPm93sj/aECK
DAkzCG+ivGYacZTUtGJz27U6KHUaTlfoe2Z6faon+YmWGIO5Gk+yz5Gh4LCrAh7qdTuoK8JyqNvK
bc7+CygQmkzRW2wZSxr1Nrv7XL4xK+FIGFCeef0LhMtXIOVwQrpCRPJqCJvJHquXZbjCT/HAHQAj
reU4I3H6/4Y6wwbnRmz3sd+aLKHKABDewpkL4VKjc8VZa3UOv08S1r0aVKERvefmnVogNrmjkUR5
DBIvhOO7mtpgNjVvj3JqIRVkGPvvePYrxnZXZnWyvdl+YawtjWJ3J+2Smz8hUU6b2WKNAJMz4YOm
5Gqdi4DNLYXJaqVKWVIJ9k8kH7j/37AjanJMvnNSY3mxxZ+3rMTBJTEX6HeSgfsTmUAfT9fXQp0E
rLlQffkHe+05wlss0bS/aZuudILHzNoqWiqVTk3yHvTX+ctoGWYwhhg5Z/t/GffZbs9q6vscCuzL
YIRGTsjLUQg8t2QkdrBfPbKIj+wn0o/rcCwscyy5wJfbC6uCiUOpTRhGT5hqKiilzKwg8xXBqmgf
UUwqHyIUGMDvKP/i8JJFKjFghK1XWxr0QvcY9YgLbiaYNppTsLKi1KRRole1Q6cFrsici4Pv7X7d
S7NiRvRgG1crQP/EV8b614utwSDjYgIf8CjLx17t8bR0fS13ljP6ndB01qsQIobATflnF/pPhd1x
HEnKgfMGkjJRi38+IvYK9RpyW/QOy6kmTWj4pM7YhvJpUlggYsvfU7RF4DnRO/CobiTkh4v/03Rt
wp8GjeVhsBErru3y3n5c/owSRiNQ6XaBS3trDRaHsBQU6l2GELkFKdAqUtqLVEofiyPUjpmXdAQ7
HcA+g1JzeruGNRC93ozhGB3fX+Evpo/GyyOrGCH0gV4Buzz/Hmx51FPOg4epcRjaxl17V+D2ChaC
gH+tIprNmc42cIrOiQUwu3rbwYRmmkxXAkToog11KpJQ9oaNQHl/GIEn1g3JMt5FIhrNB3nXalNH
T4rf3YtsuV/00oWj4GMTuHxmeASb7upWE5RfMx1yK0lJp1YctJP4Mc/YLkM6sBx3PFrlfketPs1i
svHF4hMKG2fW6F7qIh6crYOgtpXDIjgC+kBu98G9BmywBKmF7qMpQLs8Chn/igPJ77onOQCMr5QC
pmWt8B0LPcijM4CHFpRenRo+hRzJgz2kfZYSbV+p/djp51nai2Xboyvl4jG83L7DkZ2M6rMEWA/0
W8J1r+cQMPPRtDtqj3kMioFIOLhE36qcUhx44kNrRX8TQC5EXb8QcXdlBa5jfGyDhTA2IlYWTlXz
1u6HbI12G0Ex2KmWwTNLTfG04QRS1Vl6I/lz+xKP8m/Ng+DnhXTBY1blAChG3iaGTyjlydf1cy2R
sgN+XtDOEeSnQKRTtNpvAKA7KyZWoBh1KvPzuVWiOpVlbNVo9HfbAinYFjlWislYnBDg+PFXIZYB
YTMyWDLSjw9NLdv5910uiAjG+K6k8WNZrGeudn9Qvx5VPP1tCXvniOs1VSVQ23pOaj7ZCGcG748z
IZO016X37E/ajJcAJPU5ePYegl0LbayNvRIdiK35iwVjXEDj5rFdeKliWuE0BEUstCTdQhtHUrOS
fHQ4Pyaz6f9CJOBe/0nTmxxXFmcaz3jGGdZ/cefHIpGrOvDoLcpukd9rJ7WT85nY6TQmETFgpaXM
ghvWrmPNS2sYquLfLqYdeE7wKuCR2D3Uv0yQV8SAyFOtxwDfdf6aAvnufhCewX0kWP9+70cooKu2
2qQzpMhU4jBWj1GAtcrCyYBZa0US+aOfXZClruIgSug4nL4BhO1LxnvsMap3xo0rUlTTPKxAPuYG
ktfNQKkSLJ7DtP5vIlM5OAOfvQbatKJpGHHkEey2Fy8eqaxfP4sdCryNU7f2xOf9OJBavY43wF8a
+Q/iUODJDEkxef0dvSia8M+UoPH7kFfNRzFaSFjLfe3JfepfT5zW4K8pe52GItkd0OMxonxtnHHc
9QL9odqpTMobBDat/ISoO2eGR1zquSgDAt0CBk2BlOmwCC85L9zJ/ZlhLSuw3vxCypUYMHeceucv
0T1xuR6lr/82zIx7kpxuZ8iBiH+4QNlmCEDtu9/+NutqSsvP+l+RUMjA1P9TKk/k7QlcHDfvDH5+
5he5s/0BkLY6Y78OtteypuPRsYJIOGDOevs3Y0b9PYaXvUJuBG/L3FI5sn9x9BNu8gBTKMDooxpB
naqsT3VnuAVk3m09ZnLDcB01VJzEJ7PaQY8KawIM8neYp2SGMsUlMRrutQ8z/CWUqC/zjbAbQ4kE
TEWIOnfyX8SYNS0Y33v40n4iadwfVRHFNHpa/eN35ZHWQ+1FcMK01pJVQnu5Gf1rXUKrYkMV0Y52
ItDNdawPqRsuP1BGE/xkBpqSZRS+VFG807+Ydozc4OBEkEBAvmnFCCtSczKPoNq/ZG04pwePr/kQ
78ycYGbloWFho9GfhNh/i86rsNWhtl+8kRH9GbiGraCyGST5H8m2A9QmSbv9ucsND8AtwliRBkEN
kioMUPDPQblrD8i+YMkY6mcOS4+4MiafBL5q/BHqbue4SQLEX7fBwdBQoxaaFtT6K3sHnlV3Lx7I
6TxwJezITcKSlZhat+jwDufLQk03IwhwJZMo0JAQFFuJeUbpiWSQKaP6Y54oz1MR5rj4TUx0Rfds
Tr1kMVSmDhWEmYB19AUpUPmm7EFH3SYmXZ04Q1vrKJqlLwkj71SjnUeWqirf88k8qoSq0e/bYxed
oinm7UtuELCuvOGDomf91CoTRrnY6f3Vf1RI5IxN/9M0zOoKIUF/8sEeshp18N3R298riP4k9p6/
st50szAQdDnYgfvJ+rQ6WJQqS8VGF6QB/TT7XGa8uKGn5CPbGRv9OS/0C/KdrrNa2Hvw/DIfATav
t4iyAUfXQs2vUq3yr6YJdeis51LCTApW1i0+t6KCwxFcNu85bMm/VWx7Tz140NmUNyKAMhyKQukC
kRW8FIhz80a19i1PyDfQneVT2Ug00MYQ8oQPXB9rOTtehsnO0HvNYoj1lrqmmlIYyRfFdz1KU8Zx
Ea4jJka0shyczDoN0ejRO8A4DOniMOzapyJIGOhlxUBHfN7i7WLOnbVtNgpjgSlyIlCGjRD9dBG4
CpeYAJrp9pO89Nl3I2kLyPfca8nAHcW5eQHwCEFoePb/+NQjjFjqZaBrO4MS1sOqUy+GIiwliqOP
147hOEQhl0QNfQY1w/gHzKyOYvifOGgyZD6/9YPlSqeAeLSLPnGnBibaqJxhkTmNuqTRm+g6FIVw
wsplPJrpnfesfcREEX4htYKkAxnkQTMufIzxIWD1gHKmkvgkSxUVoiCzq8ooHncrPSPuLez1NqBN
Uy7qoCgsJjmsKGjZTE8ySQ1AnQhowJRT6VsFYuitw73ZGC/utgdDVxcECLVdWmbtaLpfRkcsgsKC
/te6HSfcbGrYeTCwf4DNB7neWuQm87GF3GOS2poU8mRXvfFrcMjE20AUvY/cMD2pqGPvTIRsmsTQ
tPqtD5xuSKbfDiTIiiIuRqAJJGmVRpMT5NLWphuEFNNh16+57AdCa6/IZfaE60wPQ6SS6yx7RKeQ
tGhyT53tKtkqTs6DDx0IU4rpgAeddcgNQojKKahaYUsh2kQcl7TzrcfpQEyVS+3DEndvwskK2ySU
BUFPfjwN9VZ/SV7YvB6KKy0GaWs39InwFwzWaHmWvPjdFYo66UtF8ENvjh1+lCUfp2q9jCM53Adm
O2/OVprywL5XaD9NsgelJm4hinaQ73bzVsoECs5c6mGxmaBzIe/3iejnNaKKCEpGFDEbA4SA3xnp
ySpEJXYwAvFUPk1O7p7suj4y0WZDy8VK+XBx2ZnPMMu1M2eybZ76jZx8hbVBTdWZZJpIyOlXwPxf
cOBTJ4YMkSsfzclGgnJGlfxqbgc9rKBICMxN+3pcyRAZlqf51gQpCKLgeiuNgj2T7jwB5AGoYsjV
2uCcg59uftNj0o0krRe9lYDgqMC8I1sj6ZRDXTgHK5CKILl15RvUudmBDqCX47jHMI1hzf8gtKlv
opz78RQYKONEIc2egNwCgVk2oU1sgX6stfJz1nHQl1a+M2c+tl8VIdg4LmGhE6AhWqlG7Nv7yw/0
uLINCGnxQ5Q1AWHLSKItrj+1f8EVtmXB1plvrQz8oqrVzy8+TCpR0fYCQ8u+omEcaJz9/79opYt5
SKYv3x4xFjKdSe6iSfM834rPIn3AK97ZmYafgYSLJPKOJLTPfYL5H2QxLrKVKOx1vdIDMC6qEX3R
cCNSrmufqqo/bQ73H6vsxngnTj/qxqUN6q3wmlu8/PiE8w2C2wm3sAHUtJ2OcJhVibRK/ZPHgtab
ZmBgoDd9RFcbee8+3ryvnaS5gVIp9oGAfq0mpw52HZ4rJXR5F/MFboZ3o7VGtMRNd2hy3B0PyTd/
17zVjDpu4lm4ntclpa9wuDX9Q7F+MYb+XpB7sHW1VKHRoorxVwcht2TpTYhpJAROHwzpQrREAFHF
VdFlweywnT3i08xQdyhL9bkfbdqVB4HrHQ7efLrZSmZ71r84F1IM4kffvlhiH5KXSAzCupBAmVb9
yE3E26HLhSYq9TooLxH8vKSuVMSEvE1MySTqNVYuHQs0ba+/HCaFouFTwfZXOcdSaSLeY1UZtL8R
ZeqLkE+GFMUOYzj0yyBu906gFPwhaZpvrhHRqQpRVdOx80msYijdcyw0uyOfc6Sp9bqJaYTglC0V
a9+n9N2BrBu5509sMmHl6ut/9EzNlnGyox7V9K1rssEX7jnlF5hbmzNpry+lE0e//X7E7up29uaT
NTpwR2/09wdIoqICmz4oerL+B8rsY1bTat1VtR+JNSaAaGkMaGl0J0j+H4zK+F2YYD51+ZLNQjJw
8gSNh5FWWkS6y1rFZwjRNssAMStj+v7K3AiANO9N1UffB04Qi+9vJ2EjthYkGrmBkkvDCTThsBPU
SFgwBej0tke93Z6rODfiS1F5Kxf8iCqtZAV/wIY5u6xwflS0B5Jw02IugUW+ppXg9i0haBAtfSyf
bYnIaf+uEXhflyHRtoR/x/B5sA0kRyFcSM4zpQbBsqxf42QmvN3CYntKSwmocrQVpEdFTxF2vgXq
2424+bpmGjgUjGMwpVsZrcPCCbeNLW7EwQuEzTeVlTOl0HGJTSM/KuQdsUsWtWtyGXbld+cvdu2y
CE872zxAbuu+9evaSNBXLjkdLX9Z9hMZO5od53IMLBpezQ1Y983DtO+Fe9DinSuCXenPIjgFGt2b
38phjx+q5O1lnFzgcWFEbgRSJdRDgORCRRMGg6DksYKrtaO9akqelOrraedgqg7r7u59TLuj7AlK
9k5Ns5ABytSMDf5HlVA5gKyOt4asrNw7Os1Z+Rpnl5kQr6ImiZ73SWkxD86CccEmcuFadhHlfZI1
dPaSnj+CfSkDCaj+lo0NnuiXiLys4u3/qHu10cU101hGaPR14qocQI6GXTfNmqjbUJIhEgkKmImn
1kp7Nb52BtUhl+amH9tXpHCvsJlk6v79DFosH55JJjAAooozyoYq+uyPlj/+Ey16hFgSqK0Vxz8g
Mos4MvJvbm+mtBgtU7MmYncUgK8VAN+ihn15eoIJOUayja0A3Q2ep7D7atgJTmEUf7za31pdK2ep
yKKyHJ/vruM8isct5QJuMoWV5q3NcW8y7PJub5LXmOnf2+Aflnk/7kcbFctRixXDbBROPLpvoi7d
G189fxNMjGt+Njo2g+/uSJhUvldlqXBXNAzc7U8uUBAJ7YkQfh0cEswNWR7LAcqBS4uBtMfNV3af
HnHqi8ssRL8GRWDuWdPvNr6d9cIscva5zWJetAoWU+LGD2YjOJspGf6zSKgkOft2yjs+t7IMpT9v
TszH2J2uySk+Htz3uQTWSEeDrfJD54DD1sJA05UxYIa/LmyABaFddk6YomukhYa0oMzqlQlWF0VP
xZ3Is5edTH3fnQEAY5EjO7m01Mqb2e5Rq58RrUNY7v811mpFmS3bJsdE+BIXW9qoK2kZTJalGzOd
huS3Z86WkURt08PsG1Z2k+6P45YbsZ9fmNu5GQjLfSAb+Sfxh2Qir42wVG98WEileYMHgM3QZKAa
DNAsoa5Emtx2KB7kqFguJwrpv1DExkfrM5cIunNWvz9btA8wKoyg84EhnKVlles6N2BPhwcFTh90
9WSDSJIIjqW9g+yD9sEoCmnaesNRTV8sAyTNPKCAhrAhtcTehNPZkazwnB+sUS+4QwHb3W9eSoDE
dLSpBj1QHqMAoxHJPXY2s2aY7E738PPgCaLjLLvAwzD+kDdv6/4z0h/OTgDYQWDjr0YHeqbu0k5p
IthFYt0x05+u0UNZlExEzaQsRic/+NJbFrDRElHA0E6boBSo9sI2WUz0c10J4quhAGezg6lDhoZT
p7cAoVsO5PkswxB/JR1TiwHkqBZ2Rs78TyOWcUTI1PCSciXJHnoLczZneDZ1Ah16ulT6iqjSqN+l
JgcWbw6kIjRKEAvEr+1rgWqWau9edwX70gr8NRxG0T0K8gvz+ObRIL2t+plfxhPkfL3dnkEMZKxo
2BXyYUWKob++9lHtlYvbL1XnwxuJ0aQgTwTpQuXfbT67SXor804NHi4F3rZPzPly9XWDiThitbmq
AlNCmsXyTefyRuT5gwYOxWXyhfLat+E8pukQt5dsXwG6L1dhfQgotaaY5ZKL1tWzXcRpaVC581e4
XuBEtbLA8rd8aXJE7zdt9ILUJ4DufPxTIT77XQfGYlwnxGfm4tNsHssGyaXGmLw/ZPiFL9/MVVOX
/fixMrjRzaoQwmsju2Fqx4uw9HQerGEsPW0MwbzNmLSU4Wv6fkGcCQeRMuSZBEGA6QZeLozG+lli
O2th/TGrPiuNk8kVyWfeYAcVz7wnJuX8I23+DZL5bWM+7RSEhHURpzRawCxIw9Q/xgjhMWpRVWS/
FiD/3OoZg+uz/XiMtPcRVHgdSpDlN2l/KleAYOtvrqJyeUaH7SZrXfK5mDr4JN5FLw/XVeojoTAj
mmoLL/fDAot73T1c4yoS5sC1g9xMvC6vYO1Ds2qvJoWWUsllLmWtDMGQRwxnhn/tg/sV3rQcWIwy
30I0bxDtdoXr2HKV1TJuiHsuTtqi7D3Z6PcVdYpDkoLDRE3PwNnwSfgU72FEtqV4hOI3aXUyNrnE
hOSu9nrKGrGNQI2SjcIlqu7WT+1LfA9x9Buhh2jCOVG+4W5UuSzBsu2nYHBxLUZ41Fl4vNmCk/vx
t2hf6ouSnYo6MVnNuclDMVPRLxTEe6VtYsrwQ89Te1b1WeYYa/dty6qs8wRB7xaFrny85nshRh0/
p4+dWxMPWQXE5+cKRatrpnQp5SI8C7jdpgiHxGAjk/trEH6OlRiq18n+hi1ywpMICeDytpZDoDdu
mbjqNmbkVWgYjuhPLsZ5/qGXHz9nRMvT6mhyD1YnartXJ2Fc3uw84IQEepJmnsEYnolVwVJlKsdR
At45dOcqKzv6pqAZRNpenwlAiYlGtipo8wxagJdot0TikluLq/L8QQFPU5i7Gp142qzl/8inBCvG
u1w/GDhWKywdHuQYw+5Mk1hMtm9prAjnw3CiCeONui82tVzcghGoaTbhcoi8SPydP6fqEQUJZnOq
3mABikqbL4UY+8OuJmk89+lNukaz0wTQtkpln49oQm74UyRA8amqxCLHoq/wWeUo6Fb8t1b8+zVP
5pSgUR4+ehiwufnPz1eVlBYxBqk0HrwIom/i7VoccFd4hrWsixAqH8NpvpXqCUS2xjfdA8QnY9wP
qiwq7F9DzohZfd/omHEVXWPIftFLchZeH7lCLwqZMl8aQPS5GhOz2bQ2U30wg53Hk/2+SmfRz1hD
Md8F64GGKBagqrbZNAaYKBrQoqINnUlTOVSAKLUBssihFCcFxmeghRPpt2Ipy5WEXstdJQLEylag
wV5SZtgLxhjrHbyfDzgoM39+R8XgO78bvRGJAsoy2h/z5qjTTCNfGX56lmKrGbjGhOjgMtc51kB/
7At8JSI/eql69N0kofgYt5Q5AXKv+eZhetQEM5vazt1EJ6QyBTWZsetMyJxdEVaJCA4RvmfHbxeO
v4QARVM/ggx8WlTRMRWXfKqJKIgVJe8wb0bz66RmVD8CuXfXWy6NSD+nntbbBHu5H4UM7SCPGsbm
Vvv6ZWAfOvA2BSbVNo7IdlW6n+RouUAEn+TFeE93+4aQKFgivLGRCGHp511CmYsYacg3GB276Alw
OAj7m5uCUABg22+bWiURwFGcj3+SlPe1c2DfY1GLf39JyGcPjW9YsuFsvbpHrLduZqk0864T3YNt
x1eTwPm8yiysvSLqtzWx142FBUnujXGy3IYbEyx11srb6zgag7tqoGYxKzXdSM7hG6mQflC17wDA
I4/VsvbJTi+4pP8VCyuWMM4MDUz2snSK+gcq2SGep7bytSM2WoUaqeO8DncCMD4cm3sn5yS2F7h+
byHb3PJdm5x4YHPspR7JOl0O9+cAKgp7XSsQ3z/YEgr8xbc5jf3nEG5Y/EhT3xIbYVQsPouVRp+N
PmuftjWMY2pTVS23+AgH1juuTAwaq9Yo1T0ygwu/zsCjp88RHCDPLtLTdt9RR7j8e0sp0xXFlEBr
5gEGCqTy1oihLK2NlO4uixYYlKF55qlyXAgUghaT3Pj6Mx+4aAaRzOO0AUseEOlTTUEdBxucsq8g
zpLbwTG90YZX+ZkIMxx99EgX0XGrVZh1KtYSvAYE91ozMWX6+dRvYxy/EEe6e2XGfLm4f18d5njO
qIjQ1FMHtGsIHMa/C9IJPREKSc2+JvdPFisaCqSvD36uR3V9gMsMaPAHLQTd4auHqWTljOg7JFLo
Rlq744c3BaeM1WZZX8L1nZoHBXc0H5nQasSrHFnUMNBXYI7skw/hBoYkrNNuFolxkRgFT0eiJbP4
9sv3CRT2A8VcUPbRvBe57m8bxEK8okpBdqyx5m6nk7XbikD+XVCoW/DXgPuPq7y/lIEc97dqADxv
WOUolRkJyOAV9tooHjVWvb19iYN+riLsVYSWrqiDTj4c1yRSkLzudDFuy3HwFSq4eFGrlFnunJU8
DdeT97sBJ9kdkZCdfndHtG1P6fP8E8VfSELRp5gAR+tTAoybs0Xuj+tnuYjuYsbSGGZP/uJUnhqW
1Fl9J4LivmN7oEkVxNbYz/geJ76OSPN7jtGKzD70L2QqlAthAY1nJv8pUvL8q8l/MwzGp43JT6uJ
pUz/pivMADataYIw4ju8dUIyyUf7nwNSypzXXmBYMirI96owipXSJEPeoR42UvkfXU3XzaSvcSpe
xX4nRdC1UeoJ8QgLJpO2o6zRPPglNr2aHVdIImynRICedZ2RCwzgs1YF5mSS0MABYPeRFjm1wlNM
A4CeJGp4wMAsBOn6YgsNt5oaY4gBBlTCeWUlQkIyTC5ufgJWpvCIOiHItvYWI+3AgE4D+5l123iE
sMtZ8CpA/wDAgunwzmHFyFBFRdZQcB6XWWGrlzWtYsrYqJfmuZ2cVdN4zCQRkHMXDQJdSFBGaOF0
3Efh/t7YeuXGXATEs5hKFTsy0wHgGds4HescTimiiwzNEHwxjCUtksa8WBWDsMLKzoKXNIBo5S80
SRfKm1JZUUk+wluwSk84xYtoMGOrEmQEk3Osv+IAG1QaYHpIi9XQbHjDl3hn0ru6XbSGvwJ/oArE
MV74N0ZIPxA0gINdgY2YrePguSfT9PiiDvfiQx17nls6qNaoM/IYtK1nSX1V0NMPf4TAgx/dwe+h
avn7cFyQ1yazaw9FzmWKN3vMa3OA87ly861DpgWK/+I3G++cXQ9VU7hgzlA7UndtPYpkIcuIIqtr
6C6aaYXILotcMqk28TM04YqyNVlZ491Fwq3BLupAEpSJNQ7vpFTkkt1HYZjfo16hs5bpAQMdKunZ
gNYKC/1btg09xL5dPubOXrd56fLenw0ygXZuZS8TuoLYcXZbNZociPcyHJQfr+CzQPzQXbxXAyOv
zmXTz/D0vfXWbwc5i0gYVQhkRK4lng7xIr5FBwSwSYS6umEbpqtnmxVHwZSURU1Sj7PhnXYI8zb7
HFDQmIpxa8lQEAQE0LxT3tRsoCxzbCFELkGZQfdkPk85QxhAZ1cvHRkoZITWjQ42MrsD+hseopbj
su+CgGyby3D15pneeWBi/IQWTvJlpXR+pDwNM+v6pgIlG1DLf077o4oC8KoUwNNRBoVHYV5bSRs2
EjKtlwd2tp382LGgG98F3dm5LhMnjCXcX+ZcJUq5/6iLqROiFZbvP3k3GB3rk7VGi70J6ugwU34u
OLZSsyCiNEtQRBEvDX2Mr5AIchfH1+OJvkeGaa1qKKiItBA7yNxfQE0GQog4eRosBp9canyV2gzz
/hGf/HIbc1O014GAjzzhPPiWcHPnW3u8E7M8be0hwTte/JkzUVyTdkl1BJy/avVGSDTiQF2E9YF0
HzKv1gl8fusEx1lOsZfpB7a748ELaEQ4wMAYKRXs4gvEelZxJFmDTxtcbWJHt3jP5zcRI6JXe2LW
1C5CbhgEFJ/toshaQtdOcjNywXrzxA7F2DXi2wYu2ZPuM7l+iQBVw/9JMAB4RHKonPIq7rmcHmNB
YmXjjW0hxSqu8XMtCPLX2tvG/Z9faK6IgqZhy6mmqkjxEhq2rgZCHND7zhKccINRNgnGA10pbS4L
7gRMvNs1bERM+z2pyPke6kjCBZJBlsA5UQew5/NeMuGLf+17QKd+JZY/cIWc6JpF1hQ3hyTK/KXl
7W/yO0GW2cJNqNrXHH/JvEFInF+fpgiI9/ZMdD1TmAEZjWlwAPNXre3pJHH53aaDWShOFjlJP/Cf
jFWiO2d5EB1Xs63lIg1QIYt9MjGyRMt3oqB/7IiOAXmEthXklgsZPvG+THHtT6FmHiJG2h0J57Re
ixrAxzhKkzm2oPgn2wtqa6OqbfhAPBecN+PQi5RchQWqrrFyzBPNAOPo1typ4sEA//XEcX8nzKnB
illXh2jXHxPu1iuWI2qczTFWC0YATHTKvR5PRZuSk/0ZRxApE4RMg8i3TYhpfavIvegp7BQ9MZMF
TE5Vd6GwbRMY3LZytYKRyzplhXrkVSM3sRuLvF9AUkPADkVPHacZf5z8lhFnerqZqNKqbuYTb/6u
Y7ofhLhyXNC2ixwAl1+pFA7jQl+bxzq8bPUXrtSx9ptFNtwERtekOB8xQ9En6u41WknqMXQPdANj
GTFUW43O1UFi1cjbTQFL2wVH+fDewsmI0JzoTipUD03m5S0FmrFjohxriUhBLHp6U8PCkfaYEGKA
2s89urWKxQRrNocY3o4E85bedbLkyW8JafPTW1SiifkCtfOvNgHkFSVF6RpQaWktA0bUWpmR/GQy
N0RL4TIxWwlhN4dJ7Oh0OgkdueWU0Pgsn0rAnkOtHqw6Ny8Viq0inCxO00BHhSYYXTimjC7z/oUw
qG3TiOpy3CYqoUAIIt2kmZxGnZyzJdPLNzAJ8qRdNO2878B5nd/Ys9wG7LH3bC+8R6FKt4o05w5O
jZ2CMBoaWbLpbX7oavWOdejxGuSlG1bpy6qLzQkJlXs44BhMo719sM1oc62azF8lAf4cVRneeeIL
Wg8ujfLyozDylsqlLTgOhcEBoAhldCz/5OiWffrWnSzG6laFhVX9tQGMXekHEIQ3btBL6kB5tmpx
ObAxgbL8ILKpYNpkY7JPrMMFfES8nMmxtBQhleumhX/HJUHt216yUMcRRgAdAEz5yeo/uCXPbe4t
71mtidNxl5IEcOJocBuXRDma1iVHKIsegF3kjFARrrLkN60vBgW/pAYUiJnS2qF1GJ/VgO6mDyUg
c3ZE7vlY0gxLDB06NWSHvXYluReiay7ru8/6msGh8ruqSBcL/fWIkBFYKJiYnICeXG7YR671l9F8
TDl27mJzij3cMYc0dmDK0yLnrzzgxkT4YDf27aIuW0gPEnm3+axbRUKQNIUZYjKM2Aflxc5DSdry
H4nk/HboFtYilNF1LETVD6a6VDQqBT8z6VzxHr1e9U7emssVCgVS86FRPeOv1hWzcpmO6XHA9OAh
1u5H9J1PBLX7NfatLF3LdgrYk3k8suzSGkTtM+hG43ffUXnBwyNE3S/Pc8Khtw8GJa7LZHK+0hLl
bmrpISixiXPjPKaVS9lNFWpBILY1kfD3I6ru7Jeo9ucKSyP7Z1NXIGOsmo4D72HTD/5gDs8AO3X2
mXG4ZtaW3LRp2v+Ld6K9K32APmo/GfhwF7YVkOZz8YntolT80wsSrm7TY7ovZxhJS4+RaURPoODP
IMdzTfRqSAfmtiV0xgEtfZcErqcSntcUiVUxRCfN6oLkooxi+zzbwuvU2ztvDKQzLGq4BTmcTPR9
0KQGleptAd2gsnDw3nHyDVACqol9PD/ZcVGfzNKaFeKVhuxyhpeh1ULQJgyjo7AVSj8SRfLfKB/E
7YqN/QdevOJrWJ3AsGRn7uxbWC7qpJhJeLNRpgxWEa2/pxDF5BEXfEtxvsZHJYAMNR6F+tu0AHEB
g93F/fYTWlBrKYyE9E2SdWEEpn9K/ngKXr9J6nqV/GC/2roY3UXHAYWiKrtEy2+vnWMpZtjNrLVG
AO/KEG4ioxw/rNzRHaHub6YRfo0gud4exdsthQvQ0APLdBBs1fyA4RQhMmbFaHQE6nQ9HsdQZ1TS
mhO71OVqqy18O6wfz3Leh4nzWvAPGax5oEYR35fvWRXKByqPqGrOA9iEjoqmnNh0BqiEJE2L4R+S
wadNmuVvZK6oO18c1so8XwcMo2RvsjRZ7WDX11RIcoh3g/aUZvkqvFdqyBht+1cMz7u9hoAWn6Pl
FfjLZ3/n0RELMg790lRXZhR4VdC7Rip3it1LyiZYnXbBozZjQS4AGfGfOrrYFQW4WYEDCNip1soe
jpIByNsws+l/WJMUsp5adZo8TXZvVlxc//PNo3cYO9GKMjJLTOViy6P2/2GbUp/3Pgiwa+bbrIHP
nkfj6h6CHI/DYI0CugEh7KZi8BDDy8U0LULOOeQJuPDrt1meLoudjmd9eFGdcr/PbtK0wfD64str
5yRE9UMbVaiTBC+E4oex9+WlnekL3Xef7o5FmBZT9n6JZicjvd72EYmgbZjtxTCtR397AY17LgL7
oB1tyF4ZnMWOgggmmsJRG9lwVJQrrZOET69+zQ1IGK/kJCj3DSj0e3ddHj0oI3w+E4fmexQpiOmY
VG4Tn3KI/tZZLeq8uyLJBL7KyewF32tmvXcl5agdvdQPBe/21B9lLF0L6/g74mt3nLZF092ftXGw
ptlQ4EAbfhydzHlxB4hTdgvz3AE9sRWO7oe5Hm7QasivUbHp8DKpd1FYg994Z5X7q1w0UpjEF5Wu
W3Ja6E7B8pFz/tm7k0wlsw1UAkxzEFGnvpe2THAXZJ1q9e4Ej2cYA57BxDyg9PG3KYwDyTcOogky
WYThB9+JsXJiaULTClOgU6QNAc5sK5SywaVral5JIf0qdcNRimCdn1tYY79hjd9Bmb93lYam8Kug
55kINu6xUkiRGwNdHs+rcZrLm7MhhlKjvBQ/R+V68V3v42OB0qHR/u18Vt+VgcZ3kvOgCfO561vX
jsBWkZpKjBa2GsC4NfiyyPM4NDjSYBr5bq8lar3skbrqmdhGXe4RAgIDuUKgmmoCpaedLmjAXLkl
FGlzSie90OnURXvm4qx1M0oLmnJ6/lwm7/C/skxa5qBo50ArnzWgpjmVk3+aKd7n28OHEDfLefra
jQ3RMDOCix7qHyWpBFT41D8mEyf5lsPFVYfSorUQh5Fo1hMdqzzwmuOF299LNkB0smlBe2LbbHTf
cVyEoba0/lTo5+qEvfD7TYDF+Uc2jJO3rGGNWw7CMLk7PpY+DIkXwsthRv3DlpAJRMEZk6vVMedR
p1AkDExRQhT9gWKDelWBdr/MryXywV2vR8/PrdT2WIuoOcHiFObOYEJuKIUrIPqyDq43BdKk5wKa
Us+Tt3GUeimA1un/wwVM2RKcRkKbDXxyBl8sZwTrKye1BkC+UDvhBGsMgYJ4Yk3su6sfRSCKMrIY
qAFSZhu1mdOtq97yJmc4JzOWvt+ndijhuqjgJ+ab4xHa8gVgE9Q8sWEeelvSdn8kcC3dYapPTcFK
mIh9Q+3qZzdoXzGvLhH9YRpsqS4E2oNkEZ3GHp2w1CtxoUmOzWdaMV9yf+BPF+uMQrPyR5eVTQqG
gskuZNfXnphhmBcT49QqnUWoHxJRJKVxk7g2v4lmde6quEGH/+HsalXUnqRGcCkJrF4cPVKQRO1e
jvHIKFBJlbgbwc3gsdIzgo4n4RiNsduODWhM90XU90Qx2jKO5S5VDk1dULatz8h0KWrPRBsWnCfs
AfJlgXfRt+nGVVTQBhiGsvheWb9/eUruf5YZX+nOLrbjp3H4Icgpo4gusxBm5njmzvbxSfJ/ZY0e
HmO5fE0LwdapJWRj/3fdRrAJ8MkgnJIjgLX+FhgUdrwKzJezvQ6jEe88/MY+Uur8/zyseeHUCMIq
wMWyJFBHZ9zxJVnMpRO75b++bBHePNRlQnKOImlfX2dfHkTIl4jcCD4Hj29dQccTKJr06dwktcdD
DP9j/6dDt2888ZiJVOuSnYEEhfMAXotSjBgSR57ypj4IrM9cvqxcR2aAln2SsSrT88IEqF44CVEq
+WQrflNTd5vq53SHdmmSwx6IKlAcPNDAe69pI7bANEYlAI88AbwMGgCcIc6PjiMgs0aSCE/5/nlv
nl0Bdx2n4pqBNVIozUzCcJacgzQ4FoBcmKGzSXVGPoRGTEay9tIvyvJmNhwBYFNL6FTSTEO1cDfo
conZ8/HyHN6fne/XCY/beB+xRnLN/qS8hdILn8i6jg56nBZZV7CVghqL8TcF1ghLqA5O56Ti+LTI
Tu86I+c32r1RaP0W/oOr9ju5EooRCr+EBZ7ClR3S3jUi4uCUVlhYt0ouJeVijOg/h5P9YPoreMh1
dSpl9m2D0oEDcpEcHFM0RjgcFlux3DewxZwltGV90FDZfOVggcsWZBLBe8S6iX8qLCXCMTlKTTRN
Dsx7P5SJkXhHmMzdzDVXKQK7jqE6HfGg1yjaYcTB0eQjRQoyWPOxclZcn2Xt+54lGPswk1f5LbiZ
tfeje8qG9moPeFhlA4BKSeI3RZ3hMWFROXi6Ecv3IZcM9uM1Yr67vbUYAIrJ/oCU1djdwRuwsMc7
1qbE9QP1XkMoeFPgnNn2kIXyxEF47dBGc/T1Z9f8Wk9EazGO3qF1z4jIhqLv98h7YDiE1Wv09s6w
JyvGTMNuvwg0kDMK5N/3nEOwMwFK6l0vgMyMWgPkNnVyv3E7NdE4Do53kHGylEd4XbDnbc0GbQ4r
GbczV5inpL8/vENLYXmMa5ko67m2tZLUSSyqS0ll8pXFV8nFiOJxzc9v21gguWb7SRgVQCbbXpsy
NotW1AfdjzBKGkTetZmH7RyBqtlymc8iy9CpvuHSk9qerOGAEoNthbkDoi6mbJNJYRnXN2K/fxAC
vpsCcGuO/YBlYaNF/Jz9sxCohN8amQ+ghvFEy+pdE+5z7gcHoCAPMsCiju+kH0sXfKE1yiin5Z48
1q4jWVGuAAU28h+5Rlm0601zxs7jv9Vwp24WMlfZnF4GGnpfaQKQwgSRi6nDr0nn4vPnk04vq1BW
OTNBiDqIiFUX8rojnDW6A2NufTAKUqmQ/dwAka7mAvATdpCem5xvXH5Wvqt25wYhmuLQCdtGuXy/
RwSSicUpkhFWBuIIVmKAiqqRqvSc7yaJjPXfQTbEoQgnGJMqG/5HmgnrTvZ8FHapXHNm9CIagsbN
1D2+cOt1u5ACyequMNvoj+vfEuGW4IRs3VPb0BaIg2aQnL2DtVr6KBUkh/uc3yk55uAvMU45e6F1
yoIMWiqydsREIBJyvYBbaRTlP3HiqPn4gQdcH9ydCa5VoOCoiXSOcb/r4TiCTu/hE3qvTgih89sf
DeEow5Kos3+0mexaiKwzWcsAIqhKf+g5mkKa1HhevICu5RS4jZWvtELQeI6YJGcErkKt2E2ApQVM
XEhlwb5nyypKxFY/MqDN34GXApbPlBKo6jqMTwBTHWUpgRxH0XRO0EeZSu+dRyxjVTwXqOPf4NFz
Wc1FFWmXaPno12o/dNrLgLY41J/ur1mQJ898rrcPxSZHreCVjTzATjJSmlqrOJlYe85AJ1/+ASb4
JY8+IUzwHhdPcawv1wUZ24Qv1HNvm1DyagmM6azpB3wGkcy//s09M3fj+g2kkpB+icruUYxu/3iH
GYYd1ExjzNwdXTOIjJJpbZ44UZadBXGIrJRX6Du3n6qa9Hiy6cFS4gsoIuiexOgv1oAPnISGJCm/
1uzDvq5JRGiUkdUetrrf0wB/s2/2ZvCHPXfkfUA4mwUZdKPangNOH57Zv0X7S5R5G2L2PmTyw5i2
v4fq/1PRosJtIg2k0o1YPjQKCgVDqJFBH43Ai1mHQACTN7+/Sg+UwcUu/yrJbsf0dO9JYl9UoAxh
hUlTRk0HRBoLZDRH/gdDmCpQxL8iCWbYKFrWIGAhT/y//FX6pWGAsO6aDA1jaHJ4uEBzVUgUkjFi
z4HgzPM9T6PWl8MPfQkeBJhln4bOsdFgyDXKVBIEcZy7CkOcO0S/ly3st8+gVz8w4aJsakcDr76+
TIObOT1PROK5fRnIFwVCx3XYiqTIOc4mtwY/iL73HSY+siQQfYxxeD5ituX37ot54BFvnFh3C51C
L5JISAKrSr6zkHHsFdupr/XioePWHo9VSP6L3QCr0S1Pe4bUUuIhSYPgh8aOZcTBHL9QNztjtDw9
tPNHqoUE0nVFhC53a2DnZw6/coP7+oaKKtGepUsCCFIo7tK/AQSbSbGKSxYmgFAT4eF7c1wVNLPT
TV85wChWHGg2G2u/ptmU5aGPNbm0f55133AuFnqzXPbPHS5JzRb9qjBzAktx29ivM6aX/s7kfjSe
tMOql0IogxtqApL+llMJrG8VZ6v1hK9L1LU5cvpvrR+zXE6cU0SweYFXskbbC+yzkXs17gTX2RY+
AyA1Ce72sSr7aVmYwZR0B7kQJ2imSgCsgTMj3BWAKbHZppCiWMe5ThUQCrxr653A1yf2YFjVCPzn
jpq4HRTpjIqThVJfMjuJ7YovDWNLL3BQFTyolgcCAlesA8imp0bztDke3AdUcgePl/gzjhUUXgG6
Vr6evkp0m3woLIOb+jHmY4huUIvypcAzH2XJsbGEzbZLxFDUVJt14cQJjH4KTCTLoycKK6oWmMN9
Y6gtyftViojetsYu8q0DCzJsBo1qrE64eSSaLfOcYUoVR4ejehlGHKYhVGbbXf0uUwmjqbOPANMS
kijfJdm85vuZlHBTjwJrEnE2fnmjGEKGkYkUy0fxbzyIEAidtt2ggue2JGXuOSo41QsAnGwSZC39
C0qiWB2FmnMtESCp567UZdAX8qVXM46lYrJbThK9VYY4fViRSBceDwoIAOAf7DGSDBmQQO/X4K1x
2FfZV8UPDYtue8iFdtn57R0Js5DCnrSEiuSG3CGqcwnG05E7bkKUHqw2ukpdA6ZX9thAykCpS6av
ADt3QnlqJe8Wmt4xhuPYfE7ecvdalvldHUbpcCIcyqvShm+IrBNBnmOoVSBu58soD670oOdqyw9r
VlQxlhHDed9iTUYrq6eNAv21dHHrKtorXopYNSAJKKFyiX1JQwDgrqNGjmLd/9fTnUEcHCPWfrVt
iwDmj0Iiw7CHBL1U8Qno4Yupbsb18axQQuJqAyrWr6bWSGdtxevthNPeY3LkIu+RDd510czfvtEU
epEZyenmHT+4Q4lwW6uay2UB2//Jl5cm3x3UCc+VrWHQbJ5qs48W3JIqdh0lWcbKY0reWJrFHSK6
x6c7Ofmq+gNG/rNVGafzIOAD7yXuNZhJ0iFwz4UEQGGzE49DXi6svt12r5G23HmGmT5VMi9/I/YB
fVtV0yOIKRa3F69ShuH+kNQUU7cDyt64aayV6s7+GxLAs+ZOSwV90ErQ2GfZaNo0Z4tc1zgiCaNE
5sVnSvjI0RX2V4BRsZofif0N+hK8qQ93aNH1qCISRQPHigo6hE7i2N0aT/TqLpWbb7Q1FddfWwSg
DO8/h6Nro6i950Nkn3SwgfX3ayUavQEDPSG4rfREY5ud7JZDbOFNwZgo9Ghd+6n9A7I0hBEImvx5
vLtJ0QjRdBFrmdFBfUzbXPPiO06OCpH4EqtCwm7ApRZHkReCVz5PSUdlozn/8OcIh/FOCjZaT0gC
NxbTQIHc9AxhxDJ/4V0kUsnWUMY32aVEBX7w7fPcuCH+q6gdWpoYfaJMC9ziUxm7xd7e6U00t6Ne
WrvcMcmuIfLKKvlsa91WbPEK3FrCN045UVStpZvWLjqPCcu7byG8b7iIxJIwJCiSDxrBwhAwFxFU
rU5Oasyo4YZUlckGCjPvPzC8fHa8X6h6AZzUTsmIA2qsTPQjLEseAzQlct2aCDOF6YzdvhUIfa07
kXqzx9XcG6PQV8awtYnxbWUx7jrEEKVtqVgZBEK3r3rU2SD1qshhGmenY5HR1VcyjzbKW7xohhuN
1Os2Orll+bkssD5DT+TBiw0qMPVWrwD2DHSEm7i7ROZ4zZZKhTOK65UAG37i4qS9hDVjvLORpQaY
mxNBW5x2bidBjngmUXx/ShPq89oUiEC2g1/p6s8r86qZ+QodjPND5jktn0R1AQI6KBxBmSfqwhyt
Rneb8ymCstB/UXTc+tonXlDWOerLPbgpmevjXtFPPkux6Huw4Iq8hXyFEQDCSaAEUHS96euD9wPM
lbXm+jvzsaZMOYfHcG/GsnIlPlhZ3aUYxfZi4ZjbGYBMk5x/htubkUS35yg8IJTT0zW1qlBgmS+7
QNKU3u+i17wPwDY//zilj8ib7sPSNQZESXKvvt8tWbpnVLNjNGuaZ9moiMt0Y6NGRWQOSe187gdP
jyAO+1c8ymqcaBoi+WiyUMWTvuWLSqvG0mJN3HXtcK3SA19LjdJFmjVKHVe+qoY4QSfZQdnNR/Bu
qtsmDfBUNZ6D7Fc0Oq+Eckz2Ile4/Mp2qKITcbUPT5IMmdLEAtOqb7qOHgFu+6Yp4WXNDDiXV/xv
exQUFMuMqR0uXF2HIv28/YEZ+wvXs6JnZUp/yoVo3FU6+65z2vpD05CKB8t3BqAwulklYlBD+YyE
i5os5/lo3BTHUeL0YwCunHfFdbKoBbRcbozop9IOWKqmzS8u59BYPk91W4pezJKWE0CVhixG07k9
QekZ4HCn1+laoD/hoU67wCMQhTufejnKyWFB2Erm8zuppIFZ3uVwLMo40KkPSC+XFv52YyRATwyQ
lulHO/nXIgFt7CQoDz0jSHPF24NS8fOeUwiC/SUf9Sx6XAZGpH+PnfDnIr+XtEymUmAQLKOvltIN
tAtHvo4CB0yPcfE+iOtxsVu9f9tbYm/OsSwfli6tj6vSqCGeVzmAvIBrY2mKz69Bs4n/OoApMWs6
21nGfuWwQnz6cXGedfQDPy+clZ5U5xA6zCvjOLbe/dQPeUFp7pE95lX0UWSJq76UGqE+LaRxELLw
HCmpKuykhQEp6WlvzcAx6bZ+kJuNEBpKRKiVYaH+6mkGAicYZgAlngc4buJqNGPfN+kev+6LtOmz
yKjqmUZmKInGnQPgEwrtLAtsQskKKpPXJHxfWOPFfb1dwxNMN+vxjd8DnB3eyKdIkiNkwc5zUXe7
P+HImtw0NTxp6e0HvsHW2UThafIOZKNjN4qGFYFrwl7ZsR+uMqUzYXgxEfbhBzA5qEaS4a/Txy4g
sgrnAxgC0+i2lsYFdk1w92nIEii9FQ/OAc9rvyNvzNgSHYs7lcw1Qbwvt96bVqkjF9DjMRUI5aNt
Anaciy9zY230ZY1v0TF6R/W+4f0UeUiD7ScVEfAn2B6G/213ISwgCPbzVaV0wKYhwczgkI73UjKY
N5dXd3wZ+XngWU8NeJAhvCmmonl2hky7IkMaVrPWGYOpzAdynGhzmI0tVgxPj2gHfjrJOXjmVPqQ
5H9XnKYf+sG1y55QJEnmc2IjfHIR/FBIQYUqEBzClR0Vw7rtS6STk8vokYR+G1JqFbagQdjda3ts
cbtZOWkSoO/IvwPKVFskWQhT+jbakOgdgEd5shTnRvs4QxvF9JoH13xGuuZFgEbbTqAez4yeHwuF
w6SCUZw79gQB/aYsc6inQuuKZ7WKq8o+bygt4Rus6YoS76O3oYcY0Tj6GTkv0w8TPXsud8gjORsS
2DjFnJRseNqyuraO9NUeM/Oh5QYkfrKtWRXgP9QjNlD/h2w1iq5Ku1bCOIMFQsWJ8SbT4ooyn81X
tMKoTs/I+dgE5jThBdpxGi84l3uwsGNsbzdlOWQB2pDheGdTLUQ5Zh1k3yWpJx+cWC3PGNPNMyFF
LM3OeJxxbjDbtWq25IBLBFS5p4H6IAFuetZZvHO70vC/09fFu237FusZ3oqPXWWAY6HXqEBjwkHp
6jJd+LJBq95L8LaMLdCO7k0/2dz6xODcrQfvUZxFQ9dHylIEnE8QkXVsftU4S/v/N5tA84HXr4E1
yAGFlhoUDeLldrTlPZFpvbjUj3tbVdcpGax71Zb+XCQjGBGCKgXDX1/9Y+C+1yobBpeOScf3DeSk
7bR3+RaRRsoeCoLlwvg5OR31kLwrFRol2tCaqGuJJkkSQPZcRqvfrupJd0/ZqFZCIL8YeJY+A/qI
5mKR+srUefZTsLXqNvef432k0YPIQ5NZ49p7uuGFKKeOnwtcuJYxp/Ko8Zp+mUwJ7fomZlJrPX7n
YAMaNXhhMci237YUWXFhGkl1NcKxQS1uUbJ8X2eKEepqsvNllasggpnnntNocbdhfEKpHTicHaoK
URylq9aGQYbTHzcw6i/N3QA0hxVipREFXjjccbaIOGuRv1IlbvaAxMIIXG/Fex9ks051sQFai5h3
9ieAWPUauCABP5pZkw8MMXPOE0Oyuc4bdDUZyamBfaoK0YMQfv9YI19i9zqObrYNouLTMJ8qxQZT
o+UGi3KcJMjq4YD1TOalxQ3jYWeYNA9ugK5jgqFJOeIHneYHKGE+cX/ZrRKeye+wtJbzXHkDTR3F
su159TyCfB36emzM5MQ92Wsa4wgraqCqmh/x/N+tZJpzh7CzRP0oeRAfVL5HyDqzIoaxmwcaZxde
FVUkAss8odyA58iAGJkXl5oVil9wfKeQfgu0l9NREf3RJ0WNyxBKRyEajhEXWU0Q0VpkX9vYnEv0
F6AkYbaZBKqnpF2xAB+JF/C5swI0TPFhlV/5sJkeK5CrWRjBJedgODjLOs/g/0Vew92DjbSU9Y5T
JCDjN7gi1DW/T4IaaeysvyLeTq0Qdn1U8dw2aVBmdaWoTrHfqdQLzXdixMsmwmc0io1RMjtIGrO0
1Zqaf9bB+gjkGAYfS1fBDXJeYKLBrrWiJBXJk1c0vcItueg4MkhPNOaIXg4Eu5WmFNdJoJu8bfM0
sSisBGIGMdPT9ARAzXFaCTAzaKHP37s+wgpHiNquwrPgXuqbJo4xut+16q9/Q769GsCr7zGyLSCT
mAB41LHyCl7zBlvL1Pmkm5SKuQ+ZLsUgL1vuDpFz6NyX1RRV4F0z+HHofp8uB9z2C3Ox3ewNx1OS
gVFASbxhBJaGKS4mLsIaQ4Tbe/ZrmnMWDUotXGmmodxfNDmR+XMrYRlyDOXjx3/ya0G7m91z8jzf
OzfSNPIoNhNE6dmC/rLAoREerTPrvRz2QKJDBSxncdnJB4ds5ESAmoQJ9bfhnLDHfKCySZxpbL9s
6lvKhKUZDH0DlG2W540K6u74rQSJz8ZehHINpdupm1VTTueuk2j7N+5DTBwVgyefGTGsvlUKgfpg
t5P+iMk2zOxKMyMOmldSyfDr5wNYfE9LFFzIQ+n8UeDewsHbfnSmFHsPQtyDD6tsfVgmJigv9ud2
qiEYjxaepKVfyMojFDM3sQmYAFcqxgYeP6cVzraSpx2h9ziv/0dV6M7tzYsBGOQXCtC+NEGkb8C4
UacKq7MBk2HOAcfj9eDcajDICd83x4Ksq/3yoX3w3+Wh4HrI9qQKxeR3XYcZITnSFHN/nykYlDy9
vbvxRtIpb3S8uCE1Bzrj7nDxxlRQzP8+EY5kicpw4TAg9U2iZNXOX0vyKa+L+aCKbqCBslwDNryJ
N6AdfvbC58PWMYrcMFWOxI5V+REObxywvBXSpkD5qzIkC5sog3KowMw8j0X168hlMBwz5NvaDNnQ
OaCgynlVhtUl+4gR2F1tbtcpZckCvL9qG/bS+bj8JhAidoI/uyCn+7pQ1nEpGKlBhx1qPIR/caqA
c7fYh7iBY9QUd2N7Lg9KsCjlO9Cm22lv5ET1/AQ7IlmVoFaCt3sL4rIt8RBb9YNUj8et43qSrQZS
NZTj8kaMgNY3kGhjVOCCqMyrxZO0yu0HBcBu5LDvOddqjPiiVKMFm+2L2dkKFW9me3gKqfEL+GRB
akWrIe8F2e29nLq3YlVa3M6DvCzmqF/gI73UcDBX35OIn1YbMIg+FKbgJOnzf6gzg6xM2H1VG0tX
ufSn+YGyKl2k7b3YRHQq4fgAxC7e8igHiZK8tMM6TglrAe/udBPAfFx/ae8FrkyXmqwhY7Rrbr18
/wl6rB1TDve400uuVhZOT4svWMbdQwi0LB5HwXxS37XrR7du9pBqai9xEVtQKhvr7G3WpvMVdBly
3FqBAqVJN/AMV6bEu99mhBHQtmk4NFEI0rNKMcdjY/04VUKTaxOsWlaCuOVgEZW7fny3KADRWAnw
qmqso6Ej99OASQ6sntsvttuQw2rbUS8LcsTSvC2jSUHSqXs/Hxk/mwvBpI0GZyag+NOCpLNPzG1H
D0ou9u1BmfFnBssBeCeCV2z6D4qQwxeBYPBzGLCtgPX9AHqpt2g7KafF+lAvvIBnkNVhNni7ba85
0GR5vUvx0mpn51HnlLXBpD1w2aAgBYKf96agP7RC2djHjAtUVzhGA2vjDf9tTmPnT+W2jmA/13s1
iKoR5rU7Sl7shSvIQrSlbLCQGwwSsNMdK5DsbVMWmKDv4ziLsm5xyxsyjBesJkrjwUK57kNF32+n
NNi7knuvTvIu0CBXA7u/9jbgevINTsbjucbi6/0jSPd5K4zxXuXh//Yvtqmuawz4FK/WmoghWrow
7kxQ30OAuda8S4qQovSaSyVl5q9J94mUGnP3ZXGladc2yIggbvq/9yRJfx/jjs8ZA0sqAsSxe/sQ
da5kzLtYzcvTKg9TKOqi4j9CIZbRjyv5lF/+7Kb7PjeA3ir0KhvsRJE677HjE0K+DBkSDsrj/VlK
57H9zivzjzd8hrP8rOYYUiX3x5g79cSwlfjYhmsm1J7dRZQ90utqEAW9jM2Xz6fM1VRoKThPYZu9
Zqbv9Tv3c6tZ37s3kTKdn+LAQq0jO8CoGxSTLN64AHvpRuwNf3ALWTPyNn4G63fePbgVFNOZdeW8
F6NUHu+sd4Ah0eEud9wH/iGHs+QaBbbMmb11KgapyVO9GUx569Jp/McWpP8DES0bOKG/TPNuLHbf
zp2Dg/WVh6GuD7DMtZ9HbiwfTJadRIXZToSqyyNtjdPqriM4gq3GuerYMuOhh1l6KbBWBKRJIW/z
VYEvOSw83BudMLgaoGN5dtQlCQm3+ed7klv9QsfpdzeHaIvKT+iZenO+HBWo5nEFac/gkMUiokmp
BBLjeyWuf/4TRvTFQw5hiRaq0B9QkKRjIf1JN/FTUB8LpV0WDeNkL/iUHt/NE8GjH3MDEbjv7t4G
csls5RbhKgUN/OJDy9mPv5HQymB5IgLOVpH/r24MSUtcJKJQRK2RehOzpzSNXBuAvdfVFx2yq+yo
9yiFn0pEBXkemu7qHgPidMIZtBAKylcbB+SspLOtP1bPFrsQ+Z8+Zb6oRyzBd/HvVsizWRQTzAV+
ImlVT0aok8ovcKQqMG1dz1ruIwY1qaEXhK0PFIpsHB/MNCIKCJDR8inpPibbZGdbSz1YecR52sLZ
b4l5JYFEP6i2c3SS+PmQOCIIzZgQjeMYkdqyu70XVmjGGNmL9rAPL+RDOC9qnnAG91DMETC7ztag
weQZV3AS2pRFtQoXPq4mAJfbOurfaV6GsFDNZu99N+r7ZxVjv5OEySoB/svwc/jmSVv/jc9R2Xcm
Vow7BVXgdN3stfetz7PpSqIrO1lFmky+5gR2evx8SSkQbwZhh5TDoz88KwIx3nl8CNiZE07GzBTu
Xx+6Wm6H6Ga9dilNtd5cf8c2Zg1HdHxBApJ3T3wJWVT6ArI8ZjVn2JAqCBDuLA9b9OVarinZdfIf
qu8YmmMHlLoJPc8tZhqBeLZEWyTTDUuAfuH0z0hmADS8RG5e4dmNxu2eB5j+Nw9plqllC+7WGNPu
Q5o95M2TTHThaxDQk6NfpDzavEgdqxQENIWbCGnDPypH/kvF2g4GTf8FMNjFQmv6Ehe9p/S10Dar
7ak29E4bb+ocjSz0fiyl/kLWzA0jDc3nfXl0LxrE7g3rSDqnbsPmCYvOKbbDHJx2aP/Q1sF+/hPu
ErVVmxeR+e1349SVO7ReyYioQ6El2C56Xs1f1Msus0dTKfY8kMhJQw9mObbn7zC7nZvomnmqrxlq
WwdIOoL1gkDcF9H322Io9XW31/KoyPBEJgf9To2TOcYjP9wC/za4P/H72t11GLaaHKyzGRq2Nwks
nQ8oZ6DrYJpIBPFdvFNg0QmhFufqr00Bf/j62lLTA5rZxqMfKHTgQm11rDzAF1ilkcw2w+HBAVeb
reWymcP9/cyQezS8Gss2s8NvN3pUoS7uNuZ9XNZzuIx/JgfxDkPhaSu3pbgVER4lETUA58/pN9yO
IgRZLaKjwyDSm+A0z9PQKtlxTn9VS1WO4tgsYt/YgWDO2ovoNxCJbBFlf/aMKusjT2ZEhkn0lv7S
9Rh+JuSieKv547qKLG4TZWUyUyPY91qirz3jTVzE9XqE01ECSooxUTNOrX/Y7Q7XX+uDIuEGdI1C
8yjTf6pxbw9mamC9GRgacnwR+BtMCPhO9B1txEyGA+2lGUrF0QkFtFavG61xh0BFVZ4p+NdBidPl
TJfizpGsI3q+qArgJqTXJK3d1kIpituRWV2MSCF6k/PADIFhFWNsuJiiSqRiDDDk2BSU2QqEZiYs
Ti7wIqK0Yw0A2aB5LB1tiOVzJtuT215MCAEmzmXlovo2RBpU8J+RdCRUT5bC5vycntCmIo8Gc5eR
rvZfvPWrs3iuQHb2Dru1WfV/H1K5Mo1qH+DIDbHv7qNory9Qeh5/yCYHIAQoN6UGn+OxoFUAPA/F
FJuqas8Mo02fMHgENEAwBut1i2bJlJ0CyKB4Q6GmNPxBoC6B0Vh2PVQgCOaZYkUSbnZkVBY55QAM
ThkexOZGHzH/b95H5WwItYBJqLjiRnPF+NWPHrdkLrGSNNHlH4mebbuFIfcPImlK9blZH1WYMtid
LsztNmmiFNPaq347x/wyhnL9oedzesHpQXkMr6dSt0SyeVI2+NPVvec5WNK5n+TKdvgpZvLJsdVT
RCtzq3nALM9J+L94QPPeCAyDggv7ocnLcgCUP3sA9Oi94jYhTXocBrBApeKNrMaSthcUMgIEOUYE
QTRgBlSk0rVuwJxDF+gL1WZPTJPL+SM298jWCE6umRmzMSG9QqT+7knGRnSIGob3J00RcfpTQRDc
fFFJPOazqw4d21Cc4iHBs+lc4LGjHLxIU0OO1SChhGEvtSoCYh6Ch6C23X3CB+Zk+XHAeN3/HjgZ
jIjZV0ftmqCOpCLDsTiROLh4GjPDRQNgAfbDEQF2POLdeusEnP7FF/uCYImNmp/ZTurZHITbmDiD
+4YzjPs9rKoBV6KKDEALklFqTgrn6liSZQxSvGt3V2EEORER8R6UVcGyRMBL8paTuSn9Lkauyus6
qh7mAWL7ZEFzKLz/6OmjgHuSKYHzDAxHz2geCuG7FA7Y6BLwgPaJuMWaCpHyoDd4Fvos/ZZ/bIef
LhJzYRTIUGlcYRBw895wdAeQXQL9WEa0a2v3Mb40j4VeZJXf2sPphd99jiG3KzQXnI8qVgUhB5by
mbDj+vWrPxt2wRwD2L9gXZp085vNiFbR5XOTMqbAujzCDKEN56+vwQwwctiLIMdSa7qydXIGnvzK
0gSOrIcdhT01hv2Esk76KeZJkKGEdb5yaHYJ0f4LHts7gGgjj+yrEp18hfHBb/cG1GALxxMnwchQ
BzJIaUPKcAERiY3JMbDooZhD7s0dbGGpOQGoiEj88mUL/+cGNnZp5snCBawC/WjPCohOIo8JOT8J
7MU0kEXJNIbJgUiOLOJtwU8qbYgHOq4Gkwq1RRCepMj45SVFwybdBq5cPJzwt/FMmnDuYczhk+Of
fk4F6LwSOkW0YeNyAoh8h74bEp+rhEWFqKflzVg8cfgEAj5d2zQ12Rb4ZU08a7lCoboYuRC3NDMV
udpSnZnTeaMHzO1yeq1bSG57eDbZvA2idbLCLLI6i5JA63KDnze4EvIZRf50Q7FLcRUPRT7H66i+
JmdCAYdd4WONI/xWPURRUhC1OY6GPsOBS/56gJFBGshdnQPQ/NxrR7PIS0WhTY4JgUFshjV9QKdi
YIu8ZeMQ6xR8UMD9suECYaOmBjL1hsbYVbR/A5d5hke17qx6B0OLTkvUKLFJXRG/DGkC8qDudQGd
CvHKUPPt6FX73SJYk7M57XACP0oewX+CX9nnTW1afdt7Ku48haGgPgtL5GzuVFPiZbEzCPSShx+q
wg+4aeVtdoejDJHI5Se7KLcDUct/VzV5EpYwvFYDkkM1UoDkf/hXLlt8ecbLEx9k+BqMGHWA4QvI
mJ28E1Fi2EHHTEbkppB/e7XVzncyHhM7BV0hLDwPUdMaD4ZC8bt2srKXLkrMFCZnsJXhkj7Z4THX
c3epcfQe10EFxS66N8ilHDxaFz+bIuriK54utYm9QgveECrQq10E9KTgR9avlnJ14nkobEJReBGJ
EYFLFidg5hiC0c1rMyS1PoAWLMHcciFmLRt2W+5ANHOTYUgnWda1unx+Xrj1EWt+4hiBV1c0Xt7m
Ln7O3TBEMSuY3AYjlBMC0nceip22SAIlRk8no2mcxqKEV+R5JwQXoaH00ZYulxZYOtXtQp+J+RsL
+D0WvjzzGX0unqf3hK2LTukrdHdIXUH/04+GCHgd6lAmjOOVVSwHSKYJyf1NFJFaWql66i+ih9g3
MS/D43Ig10yNQV3W3T71Cj43QyTt6QPiaeGrHbX3SYqU8hQtCJB+W0A3UW2Ds9vgim0tUWCC8S8H
crstHtom76f/iHEsDE2FwfQ3RV/M4bLCT8Y/KTKax1agEPqgpUJlJgl+2uixNCo04LmimwKYJXGq
GHORx9fvh9eEVTmyXcWmwjde6w9CQGuy24ybnWqoou6KH2RnJyotIu1lejTKhBHdzzh/H5ADS6u7
DBRCmR2IZHoiXEQjxAAjCFWfT5/LLhZBBmx4DTGMGKG4qb6hkgFg/CDFA080hjPkZZtSV0mXPFJR
JyEDF/WZtRq4oTutPJKtvRyBU3XZeob15Kfe+gEmtz5U6OwL8RgDmo1FVZBD+6/rGYdVKEFts9jz
rtrU0twnq69M7Cmy9oAAovWlH87DhoWJlScM9J1HxMYkhgxX5OS7tY47t/9R0ub2BZ9rMnr90eRj
VcZnO+1hekcthQ/3DKYyOBOclzHj3WX75kj6dl8J5kzoWMmkN9hZd4vuOrml2BotlV6xs7B5YCa6
mXnXy5a3pZsrmfSBTykiicL7xWSSRxmU/UjimXHio8UCQCom5NC0wDOSNnX3xpUmlH+6+O5/XJsL
ivyTZVmPUYjJazQAmKBZ7BCmoMcpGxvHf6RqADS4qM6Rt1ecExOmXnBZ3SSqWIboIBL3Et3eQA2M
nck30n1NCRSEWDhrXwbhD1os/4spwzdlprOnZclspU2sq1/pB6KUEH5j6iJm0pPP6rZ/3b9sz+6i
Ph8eiMPrICx/rUXKia6w1GE1XIrVDiR8h9mMvsQtNLGE8Ikq9Lms4lmEgifhADQoX9SrIZTADym5
1nN0aEPOPrk0Ao+o81BRto3qtX3C8GkMp1KXxeIGK6eHaGUEQfb1v4qSbem+KvUsRFyRUlCMYZ1R
6OqWW9gouamGxjRzJOQdHHESvAIZuCEDF4q32I/2E2lHlqi/hotBMl8Nu12YayfBDoEgxiaclxrP
pwKk7Wtfv7RrPdlsojNtIGCwCip//vBwGoP8r4AbM7qUHpqAI6N4rYxGiNagr0olpmkRFJNNjR9W
nobFTSSPjQOHqafYtYVvERS8agkCz7XOzH8qWfyX5PXWxhhOOCrxBbwqw8QhutxMA3DiDWb3rdbY
etlpMKcXBwMu+PF8pQ82bly9bfymw0ub9KV6p4MeIiV51NdNbyB6MbdiJUJ/F3BBh/hDQnAHNJWY
MDA4Y3nWVZb9jRS9M6keqCC6sRtn8OaWj3gUiJHLXY2kGGdENJ1VGLOLiHtwiGnrZJudR+P48Xoq
dEer3wjvgnVcZUFSp1FBUC07k1PJo31oE0W2IpZxIqNus5WpacED5GFYWIzEjiEqJWERyYgaT+Mw
htEqrPqmQYaO5clbn+XPkm5S1DiFttLMadkEYo/5MAR6l52lS9G1QNhvIBeqgmkwKhtGC1lqc3Od
MOQO35ozpQN8zwQ7GOLRzDjWexzVIs8VlZmxLSgTj0zwiDZP5D4KT82fE05XTq6b/4vFa1dc4XuI
eXy98MlpWvpiX0ctpRUUgCrBn0JWHMIHhIP0O5ssVnc+ZwCzXpSzS2ASYSrzDTmH3Vf6mK5vo9mU
FFGNHWBZyfTCDk5jsjyaLRx4zreVpYtEpNuYZzkEO2++buxoJ0ujkv3SNNn9jSKRfEmB8U6BwNVW
JHyS6WdrIiWmIfw8Rw668TkVS25arXLoYE7rxLw8iPbL7D0j9bOEKKdwVuw/vnyTLglOPA1oZMtt
EzO50ekpZM9aeawu0Pnf8MpfHpq1uePwzrJlcx1WdQd2VxThP7rN2AtW5pd5B8XG9YWroqmS2p3g
SAgAAJF7Ssk3NvhuBRw5tit6kKeuQ4eLzqFJCR9Jn9hAoc0vU8e67RXrAa2LO1C/Ig2lMhGqr14K
iTG4F2mHSXCNbh89DZ2SdHDlBy5fUx5BvnkHxyEZCXU5K0rPVqfDYJ8KwolYAZSlCIJ7omR4NG9a
I2eW3cScXrfjXdcgNkJS95Y/iQRxSrB5IOWb8f687LnnHEAb2zmg3EXDFde+3oVvcYaBrUtDjMoU
aqJIgudZe++hn9t4WNgAI1yIfm7QP64Ix2pZjZmXmY7005ANV4OmY/SAPBVWDOgljQRvCNH/z9Tu
6X9QQoNckeHHay+dMEmG0XaSbIBEwiM6l0UoZXt6+JiTQPquDYzi6394/qd06d333QgCu+MLsEGf
KmU38k1/pFgUZjiubFXeL8QypTpW1JDFvPfu5OwJsOG2k37xyACKG9RZqNup3OQikXgoiuudQdOH
tDiAWfGTRBkz+HoVtFQPaHUH8BiVOLnIdfG4NM733f3mrAOQ5BH3KzqHNG0jvjBqMJhvION3HBCO
BE9yEjLuAaAMtpPALeQE5BxMvDXelReZasVptaSlSCSDt9mAAKnZ7vAQ6Ga1zE5PNkA6AmiY1q0Q
j/52rfDoMHDdB6M25UnmSCEEXNtxSHasfIl4xP+46gg16tkVqlH0oGnHxz2UbsBUhV8bSvDsTy9J
Qt7WKF8YFK1WbGP1L4TFPXJTQ9MjeFoukVp/L6GCgezo5Gr1pgD9BaMmyYZg0pSfbzQUw+POE750
ImXA45uNKXZ2vlT1sTtjoiGT0ANRSm0WRLFUpEXIvmJX3wssXIiOIpjklFZvfCLR3l8bw8KKcrGY
erpIiJYPyCS7iM1VO8Wcq3yUqukDTKfP8DiAyk5gjuo3XWsh2YuCTz7+pzgDagV/r2oaXt6iaHyP
EpiDgkExb+h0f5yXOk4+nYMKKLltBOMDEjQqHhTDbRQq7n1ghShVTPNCIWU0GVwlAni7QwHUrIx5
i39Y/tFdP4FZuzteuYTZPlaFttJTB6gloQKEsv1lkhtCUifvlUSpnf6fqTGgDDcPiCQmLK2V4BZ+
sMYDlKuglHF2I38/QZwrvsyDBq0nn/dU/BPdbrupB4S54IwpxzjGnXwiH2vNLIPg0ka2pMLUEyTR
J0cG8RC62lUTQ6PALBUMl+O9gKuSjWCvitwrYvD/7nKvnjgtwaFcnpzlBhvgNH90bEWQfSnip7ql
gOFPUEyU+HF04hZL2PjL6KMKYdkdCn5qg9xnh28iwoWBKzD5izjzSoc15R9lOfyZWQkn5EWdSdYA
4tdFral97MwvygQc9/+Oc0dXNsl5Jqz51wG57LuCbLhsjHvGOyZ1OV8D1Z3j0ZrsINf/3FPb7vSb
C2TQWYDhnh1mbPElA9wAiNMKPglEgcC49j6NFTsdJntw0UUiabEtcb1WnlT/ka2imoIOArTKRNtj
x0qAGWW9qrwmHLULdWfwweloEHd3DlDKnyUs9/XX7KhGCBFc4WUs/b2AN3HUaWd9+zW/Ew4f8pQ7
7qEbJYRfBZkJAKJTAgvVx6UxizSrp3wuZiZ6E2pgo3y2CC2Pz2ujCTvkBlx3VqO1jAHDLvB3ymyk
MXdTYaVHSd6IuIGtGmU5WN8//pnui2X1CCLm6gEv4Qn3b6RG4D7e5+2lp4AKlQ+AB+BlQyzEIAib
M1jaNQQckVtFzLugB4msJT/TqpNfs3iYkW3Lsx+igWrdQ5eZZcTGGwd53J8TXxQ7RZhIxrNWmz2l
+XwMGik6D2eZd07tRNoXxLYxwIAzV4qxXj13L2dpwrkEqxF7Y6Gbg7gsFCsq3WtmMz8mMI2JOeRo
DfRGZQklmNS/6w4l19BuuRHX0kYBQ/x7dHXzpcaiNNZGLMTfJtqj56/oVbQoOP+tFbUCAHQ6cjud
2iUqpwjA+uNCjrEYzgrP8LZbc7Tz4ekU8uSY1UBHNyMy0LVpdLg6GAe7C0EqGTEaarX8C80rgbsM
vO14DO2Dkh5afZ/V3cI3zQZTsTdX1z1aEJNUQ7PAl4c23ONFwLiu9CXNeyiP24GST3x+udT48Q2y
fSCjhU2U2NkFqfqWojdldfE5CY732OuQz0DHAY2RXzJhg9yklFVOSCD8d4nWkuAKgzdCkPEoGA2e
HXgpZVlzu8qyjVtdZ4IXHQuzMD5JR9WBZcjTzYniH11b1ilKIbbqP+CcEdpZl+xM4+ioh2uzS634
ERf+pDtZgwLdcXrRC5pcPfGKfi5QNREjYDZ/C2GMTw4dFNTbHe5ehze5ltnKfMQB4b3riWUYKjhs
KLE3AqXeT4HovuQ29ZVaAJ5x/dvXV/ZHCSoXvZmPhPhg54tu7ApL+sqAuF+SHYap2l7qNppuP2TJ
pCp02cY3HG2JcIuFely7w/tUYpCIr5l39n4K+nhQo16uUfZieMzp++YKn0fSQgVdhCeswsh+xiTF
G793nU3xCcXVMKpKDkudntzqdrzxFzMYXXLOw4LMDgip9tEZ9UkFjSXYuNRYPIgby/rXqUbxypBy
rraask1UE3q/4w5dWNTIX144Lxijb9Sut+Ityyc0Qps1YUbBe5bZsU82Jxsh7IprmBQsGRLJN2rw
Uci4lvtQ5JRMHOgG7zcneLy93WQwtw6vErivoUp40hGW0/VOweb2tZ+BXk/3Cd/4sQ/kxfdCjaCm
6xIRD59X4Bziuvm143jM0lULcwfSuY3YB/Va2yN6ir8ljDJJm6hnuEk/Jhyq7cMZhg/HT+1S20g0
vgDNxfdbqNdzsI+1qAt7j92BlgBWGYsJRHtRYqL6LdWrcZx/hTHH7EqfxUMEeyYPpMFhUxxMqHEf
a2hDUsqdMTmwfqZKI6a2Wfk0pav3MXx0tiNE6iiZ0zgcNKtZ3y8UPKnL9OFA08+NIwS1N+EsEN9a
y57uV9wnBz91Cblyd5QXNbTU8ufcKqgvfbaUE+0ckv/c9pdYAdA0SjmpLVjsOq4I/CjD3OZfkH+T
Lmj/64LJ8P/JRV2AWHXk209AhZ2RYD0S5QkAiCNT/Y8qZdswbybVS0fggwDwq8tl4YfrgkPyFejq
/cno/zrEVSZOC+sBsg+laMv52y1VckDWgzRA9cGJB01Q3ApN9WcfuUshoayvvHcqwul16eT+9KDs
GSoiHZkcqizbJmquQWOPG4GOmZeV08imsmp9fYciWLZT+0Q9BNc9OEoCwzhZf1OpClYWZYvH51fc
KnIsMO+ZUd/uxVR9suBVZ+hP+G0btCEXCp1L96d9TU6ZaTAbiUG+Y0Nfw8zLVPuhiDv5VqMvR7XU
6Jt0lfJVddoOQGBRWkdt/WV2hWBvZG+id98Gb8KH+86cdVysBjFM35LvS/oN+eJI/ltZ5hCQY4G3
rLXtBAWf9aqZ41J93tSCSmnGXBHMHAZ/b785r+aJ7tf42meeIRYixh8oAvFZZSHXbBL8N+pfQDgi
kuXdsqm/w/WsQuENSjazQw++5GrJHyPDmZ3yDerpzfp/ym8zFf3GoaDW/0gWI10YudkQfZy5XrD0
OdGzUqdNjPhCQJ2ho1jPMWIQYMofjQd7Akc5pjKk2zduClGW3HFnDGeNXto2h2Fvf62nLjxpCiWI
Psi/xFVQmGbaKWfPvbM8DJjilt3739/xlMBgLwx/yF8f/9dDvyz3pD2CPGeLfChZaZKaq6Mix3C5
TTs2IFy+b9A1lZmXDiGQyXSuLNLzTRyIpVAbiSha9Vp7YY7hJ0D168A/yHUvaE+haaHMnb94Fexw
49uwAFvlU/PtCDX7I5HoKHFshZs0DMyrjvm9U6Mk2mgpu8qJp9DQCHXOXyzZQkDrss1eBUtbxbB7
PQ0Rl1Cg+pIoClf81ac+3tUVAXc9MsUdwCsTE+rKWzHqlA/C/r+saunOqljyePpeQd8ckwRe+ap5
syx4bBpkphgYfmsrP3+S/nJM05gmRgXWA290eEYdCwGKBrS0sXo73kDN/8t3Xe3Bc3nAhZ5le5bP
pvD80OL2rSxRJUFvwqqCY0tCPxtGVdKIlv//dAMRoOdLUIDB32UEE+6vlFB3iGKC4QDXH60j/h3W
f6dpnN8RpsMs4tzve+C6gTYmPMbRKKyrotb2nFv4eypeAtHXyf6QxvhOGHzmQib/g7Fiaiu0PgGe
8qlohOig3QZlGrJiGqnDg0xfz3Mkr1PpJM+Q0GdSsujiQYJNZO5qncpYIAkjGKpvFNTkaFxlGoLh
ox019uP1jA4z/De8E+Ckyq3uwyFH9omwqaqmvoZFtyofT8pWdyTPHpZ7x3rmyXXEmU1JBDrD/o7j
NPohrMJIbmUXLSiVsRUfEMuRuIfG9/1tM+GpLxvExBrygfTL0SFZ0wxSYVQZacGgIFBgzM4R429V
IzZFZCMnYQwUuRaK87Og1OzfKrMmIikiNgEv0AFcI1DasX9pmP9ginrz+RfqgTEzrax/u771szhP
OnQB2hWEsi8jQTeJzUHLx4kWk/FoWEZ2cMRnAvi/6KzZ9z8V50yxaClCLGFs6GWaXYX0vKB68J9E
yJl/Fpa7WrV0YrSBzWC8i8zRx7GQVDBNcupRNYauooYXeJwVDAFSDSFi0ygOAIUmJqIA6bID1rkx
7DyOv4aIKlDunG2fARUi6wcStVXmkFLY8A3n4qrrq27bmw8zjlT9B5TLyLPagVog2ESB35+0pcIR
BVni9c0FRNnWS5g7ESB5MW9UrqfqzG8A0Galy4wsUMMd3Q1Be5bT7XC4i3rC0Ddd1/YdIeRWVr7O
uZr0kzFfyYV4XRzWd5MWqub80mvhQLIT50AadiPJwqLRv7TbXcpr9zhV9OfJH3WRo+cH9XU6NduL
ANQHn+JICtylyOt/PzDrjb3nsC08kIY9e7m1e4tOB2iiQ6j6YbeK6bpyD4aiUBhF71p1RNebikkj
sZJOexJwO7/lXIF5q8h16M/4zIyr8Zk0M0nj0Z743py2uW52mWhLD6JpaCrrXN8Gp+Imact+5jKw
mz60u/zn2rUmSkTTvxh+UJKOXh1BlXXJPi3bdVKgyTEupwyUoekgJLXJtvnPU12BSvKgELz/YGnu
viwzXSf0lBk7fELPvP6t1r+69y/WIe65zCoYDvMKX5nKTR4jiHobvhjq4UO12DGpDMJ1muAdb34b
ga/Qpxn6i/ZwtFm4W9ysM4qPbxqLS2diJPAG5m+iEmXtmuclmxHAUUWA7GfXiwkDp82uQ3+SF94y
5iOXHN8/1Er34YSu4O5yD8nDiNH2T1DSM6ftStWX4bRdrwr87wjsnuMuxGJ+dLEkwSzaaxfo1/Zr
yav20mcU752d5mxSN5xjoWQgaVf9Z4SY2BvGO9yEAJgDFK/KWmry9YNFpm926ZjprUEwioDQ6/Rw
0J/chOUgKVzBs4vmCDaNLHuBNBmviDw9S9SJFbPRuqGujIm1bwYmYWF0eaK1q6jmHH1PUZh3PFdK
Ywf0+ie7OM16oD/sSrT7PX6SY8aRvCgB+Ztuf8zupOCXWZwfCOFLqJTA2cacMALeiy0ScvGe8uUZ
8kKXRwnxdMxo84+rNeVttrAmPrw8uNFeJdHSRNTgefJuVzE704ruJ80r/uPirFRLu0sLjoxIAaWu
lpzMndKbXDjCHbyQlUVBX2MdEWiTbdduiYkM4JYWe5ADh4HeawD0XoEietschEzBT3XZPZmYkCXl
sKPViXMmiGpzg2i7WJ9x9kra5XLPuHDBXM7WE1P4nUkR69oq65R7XAeLjFRyYv7MEN5kchu1h0PD
UDbpJSkOUMU38yAZKqvRS5N6SnQBHQZLq94vPKOYJhooK+HhvBd6aDF8jtFxS/IR/DTCS6/7429j
nw7XHwrMvXCs250G8sSJKicP0GLug/BcluURH13ipOVREaEVDR7JjD2YMy+BoB076iJdWlIkcSlS
xxqo6Mx0fZ6pOkzMr+wkxI+r3rn6hKsLn5OUix/f6puP59vmzuVtdsKbGmTHGyOhSQ5mjdd72C99
wSP5EGWGRYXRxsxXQSggTQRr5xzrNdy29nDpDIyPvX5q9Sv9VPXWIYSl7YpLsQchd4uOeiyNUEkC
L2WofBkkUJJuZDuv33ANUeExuENhmWEzcw2e8FRoc9/+OeDkOflRbsJNGSU+TsYoo14P+kjdYPHE
OhvtAXKl7+6LFwcus855xdbRMn/mZJDU6hfyc5fTP/ZUVAOtsFg3wLtjFC5k1Eu33NcQVU2QWoyt
hItSaYpWZbzgjpK5zh8OEUR3Xrs0oq6DAufjrJQ3XZwiA3k3uG8pYYRsZNxUAeKx0T3I/Hr93LUN
//o9G3QyQzfEP7xoSajWY6JmUzSeMSj27VUkbV6F8P7TcED9+hvo3p94Kpa1Mc79ftyb9NVpzfVu
pWaEd/NQIDCp22v7F+vJnqfLHVaOCELmFei00lJKvLXqBbSJmPLTbjwXM7HXz6c630T9do3i37wz
1c39jk2jVsY/sHPP7wO9iYaLyTtiNQU0bDixlMDPMfPsUpAOhVh+uyzfK02cS9re0rBsIHGT5jGd
X0eJv9KuFT/X8FtQgBIcfN5XL5ft3lKG0huN0Vkslsu69n612TKZexfN2uZ/o8DSHYNVnB82lV5+
1ZIs+xD2wBBgXPTrkPlzzu/iHqqunXtgRHrA9CXJ47UyP376KRPkqABm7+VNIyHVP6sZQ2m23bGC
B+vbIiUZ2xeG3oYJUephJJXOOBQiRQj12UrkIzPTAVA8qXgExmm1HWonrCiAn6NB5Nbnevzy+RXR
fN+xQdZDVHrV14awUL2X6wsc1HZCZhmd1lQvvYKzz7PVyhs6Y0Ta+I8fO8N9T5cbY4xk5b5Zn8ii
EgSEQdWTnAAAadntqjI+jQylsfdDwpt8ssJVZNlbpKkeR4bIbODOOKbBAr2mroE1E26OEKAAT79x
kxtJOCbqkO0+4Vzvqa+WXk/YnmDGRCeR8YQgglf4OTzCd0EGSFPCBUfvx/Wa2n3+oJ3Ihz6KcjTF
6FmxJb+klV57bYsrzCTH67m5SgInGW5gKWt1EXZVgXstgfJHGbU6D/69YIMMV67xB4qhOY5hReQP
u4sf2wtO7hkfZh7c3mkZXjT+wLgoyD/zYNd/qAO14UEH6hC70RYDcTkEp97n0p5x+l+FHPSYOhlT
TkX9ULXCit6WXDo8cMVfgQh7T2bPMqFsq1XuB+EaqTClAh4/nEoOB+MB/0Fs9fDPg/qBwX9u1KZj
Of6TXVy18rU4+nh3mR1PjG7pIx7D4bFiFILCiJn/KuXwcfGBhtdi4Zsa5vtuqzy8RSrqeiiCKRKC
ZIHkHw+LU0XLDjYoPEnzdf5hUkiUq3/uMB5AE3ZRMpf1LpBPV5awKI9IzvoA36k5MvSBX1Q6glSY
cXAIQdR4m5vYqpvmhnx5Uw2W0iDVqbONKhh89AzJAwwtSd/c+3txfe4ogrbZvf//xzQ3izxx7gZi
gIVE05aOGDsMZlalERlH2VC6CTp++/+MtqsfkgqAoHfqSUT7hFRseeV2nlJAzNF6jRdJYHaMJ8su
orYBqq7XLHB6kK40aP1PfssXp04rHZ23CSMurTwvDHquoO+IrmlYouow0mqbmmWw25XFLnJjWZHI
K6BiXCWd5kHLHd1CWJTiMwWLo+AmiMgC31xdFEEB4gUadytpRRs1/n0EQA17kw89xOHBfZEpwosX
iFVA525Om/UZZJ4McqksIY2IIKztZj9ItsYqMb1mOsf5K4aIMQRzj+/bYkEq8JPiVAhL1LtvShAj
MTACoCPeTJSpt52EPHMxmi1Ny69b//BwwoCn/NkZ4OQ6l9IrjxW4T/lW5Ua4AUiFkzMziID5xjTz
4X0fNkwTyS75mqTLlLSJdaxCeHH9pn9YGMurDqOvnfCEH/h67a4y1Wd23CrFIn58GYK+FU9BP6Mb
Mr/kyrpqa9xkMXHnHmEBp+9ln4E6Jlz2eVx8npzYi5T2zqT0h7FTDPw3zHxNO6OUbEqu4Eryp0n3
yhYmj/S4jPNKH3sTeE4m8fuLtmDojdsDYUUik+5IubySfqfVvLgMGMbVHEMqZuE6/jpCUSwi0TM9
vomjbdLxPNs7etrYjCoWSjqJzMS5C+YPx4pdpGkTPEC0rutzbWgOiS53C1WtZqKBY95R+t6+qKmE
7KvZwat3yT1T/hp6tvQyMDVzYckNeOvVnopK02f204fAa4gz73qu1/8Qumwzykf3miaCNEPYtNOp
zwk//2C5tmei1NJL6sVTWUEFVMu6Nj7CVEQTBrbRVKlx22oUPSRAf/tPIxeFqhxrLditZN0SXSAu
5gbqDO8xGOhCe2axTJi8SNqY2JuUFweFjaNGQW6hwvwiSD2qSaFTcKQeJbBLUpYG1ulZGBNFDFKA
cH6uWz5vDiVWGl+SWdtcmcgigYXo9CZIgTOo8GnckqH4gqL507O3OThwR32e0ItfjKYp8+7krSxu
bHhaZkolyGEQDYeKlGbFw5OpDPnzqeDzTREwiUdkqN3/0aTwuTEiwAA5mH5ILYyViOsKL1+nHGSg
Htf6qpe4xopqYClx64/UbqOQN1TyBGpUoJQOWdHiokPP91xW7FyMcVHgsoNIFNnadDUu+UJwm0Vx
G2wU0vNQPK8/uvDBYDsyezL5obeR+04HHbk0IbVu6Ydnzu3tx76D49Koh9bljEvkx1FN0YzbSmwP
/zU/+4Pvlh4cbljO6IUK4GTw2w97lLLkxd0SB+gD5nRBWHINYoKPZCucZwEpinirPbp54RBWALWd
yjD55fTj59tTS1VB7K5LwYMEIkmiSLXeLleAWnYPR2xpK8kJRUEP8+Xb+/Egjig9fYfQ2eFPFWCy
FbxPfbZFS/IU9QqbdN8hJmKJzhQ7+p1syOcHrfDiRNUnO+oLY7t/CkKUGbzMTEbugD8Xorq5W1QU
xmCZsITPuHRv+ckWNe1tjUrWiAra80XHKKTLrbaHTxw/T9BkyHIqmZuQDpgxP5H70r/OOjNvE5mb
lDni+g9v/gH9bY+qjQRH2n6JimwWcC2nq0Jswprh3hR0r2D0UoYQQZ+wLhOUZs3jorRggO9GlIxd
z7U7rWwtu30Bve7z0elBJ/qttxsIftUBfCoPhmtaPf0HjeyBOQakt2988dKYFEUxzwKT+ALOj1sr
elXqYDpQ3+fyreathyskuKzwz+UWL+IsvOq6P9lgaWWrRcuj7PZUs26U8sUMXLXNt9sRQumzH3iC
1BM6SeyIFDI0eUmGUmLxtt22at27P9uP3CUMBmZ4IycgS7gNU5XThXJufTx+QXoN4/t4/UHiJrZc
xuAatVkx8NqHmi0WKOKME5OKUWZs3rIJVgOwnz06FeE17qNhVW15hxNWZvje+10rC0hJFer+CXHh
1icY8ZV7RzFkpuSqve/fcmTqdp0Y7Tw90OSnEoIYqblU/NhHGxLzjqSpGNh5jTxCurBl/1befQoC
y/Q6o9RXrTSv3INBeYBpiN7tPgg5M05sS7nTm9t+fRJBv8xKHV4Wv1f4BBxIJrHEtrZjMmAWvJEs
N7O9jUT5BiYoUuViyRbNhFB2wstHWVIRee4tdky9S7P1P0uibJ+O0CTYf+oxeZiulMYc3DUMkQuH
ftT29tmBG0aMEbBojngFtBeEQ1jiJjdityZ1PWfPCKKgiYAZHfvp3tp6fZPuoDWNlWQQvFus5BZN
7CwcgNI69cuJhpq2ufjKeNEEWOZs2d82LfucaHL1z3XhVzykZehEVtkaUORLGCf1UIRkKG/RwPKf
YwN0Y0qr+nRLpe3RwyNa1WB5dXSW82H3DLPpS81S1x4dJooruWgGyoAftzlQrAIcX+P3SDjTm0cf
aqLRwN84ckfciwP2X3VY9ug5VVVCo4vQkkZeoV39fxRlXU6QWgO508Fmd4bxgpcs6DkrcPpyHYrQ
ragisbKzaDiEMWs3tokhCM10y5SC/GJ9auCh8r+hyIk/DtYWVOXxs6fNOrp22lQjKFDD3xewTYpK
gfWJLC7c8GUJfeIqoNLXUW/kBDxw1gvpGzntjfKNoXUSafDDEnqYohcel8wcj7b5iI5dg94Ozolx
HshKj3SL16kc/ABOx2/C0vGGX2N7rB0/qKLrz6u8luHaOR8MhZOdhuhBaXf+Vg0KpW8MrX6Y1z7G
h1itQNm2OVXUZ/RPFPU24/xsAc4bLsertGHXUNWqY70Cc5nfOSTaIIOGFVWyrlSHUPmqwSIzX4jP
acy7LwFT+O17DGvceK+z4izoV805MkVvUEv4gB7PXRs1SDPNWmrJnLNO2q3RuLQl+8olbZhZcbFz
ySnDNMX8BY1d7e676W6vCPaBSbIvpHP0JpudEpppNSFnuzNMKw/EX9ED76VCDVgyrdpsmFAzgnoq
17f7GrJVXVRqh2qMmRTcIUolVwdfyyZ8L1vsowo78WHnKNA3Y+pDaNMAWrRzKdfJiRO43tQwDw87
tddQYG/oGKkOChg7/GfQFKWaWW7YeKLqmqGlvVxCM121x4K6/qLyyRjfSrMAZ4LtdCCakHVw4Nuj
gNExJpJs9K+kNzErgOPkRvlol9xykpkXMBWL9LwSLHAeXYEvKwqiDh08XvbPjJbWmugcFYy0SjCf
ANT3xCp7fWka9ppt4DAqY7UgMeD24fjZK7pjXfhcUoBEHcnrR4HNqGwU5i5vMIYnVYqdFcRm2m2+
DgB7w+BSp7jbCF9j0uiwa8oL2tGiskrT6LxbAsosEJRsY4WJujrcYskIgkqJWKH9GGSyU/tdzsNe
+Oxo8f2UvIJTi/wzFQsrrcGCER4t2nkqTVLtrbb7kxy1D0JFt3eqcycp95+azAMJwawFxjT2R0mw
6jsngACpjM7puoMZ/t4GEz/6abZJZPARFYlsZot8ChvaCayENT7msWpEZVpQS2JthHFeXnUEkpQ7
r+fc8JpgJM6XF6WXNtLMmQawyvdWJuoUIChIWJwiKhHC29gZscZbDPuZ8UGSH49O5t2fa2hGnxOd
kLG5ehAhSQyQMMZ89oPyocqimtO0mZMo/VhO0xb4dUJkIsgHrBPmC4ybblKEHCOCxdCwmLpglpvi
dJUDDhhx1rnhUapv8SjOh7eTwtviDsW/76Q3PUDD1aRSu+1DS8WEGQh56KWNnvmknZIKSarFB7ez
bhIr4+N3PaScLp+OlhlGkV66bp7JVZ/0uz0ghYu+Krv8RqDNx4ReHCz05ROjdTDzBB1rbEmBf+e+
pVRlwf4xIDlMvIxLwm4BJH7471PlVPBVzZ1rXeWqpfRA/KPiShfPoVyVbg+9go8IayQoq1GA0yKb
BhcXNnyQ2HxCn2fjzzbJaojR2EyMxKF11xu0Shxx+nQVE3ejUIYxYFm/g9f6uQ55ROH7lqzjYpuq
QIzLlfvcad989lCblWOx+9ng3tfb5bJssxqIcMndokDvnaf5hiBqVjvibQRgR/lrSOrAxHSGDAVO
veUOAW4PZAZ59OSe/HtpmJH1OrAlk6O/9Bsk20HPJFVEuqyIrnEho7+ya9TkbW5ysCu8k7B5Xqzm
NzBYIzYHoRAFx1ni4Lszn8uCQqp02Ps0wfGUjyGlKz+jRwdtqEMbqv0TtLUm7CjK7DTNYjN3e32C
PamhTvquJmYtM5Vxc5ZeEol1EVO+pa6wTQbxzHlX5rh0h3IFWVQFjm9LVG0kQnjLGD5u+wdcEyON
P1CI+xAPoIUTVA3PnhQAQMuX82NRc+YkXrFwnqslreElFTD8mjFA6SofbGgtIZCn9sPKobJblzfU
lJw8NLoROBUh7wf23cogJjNtisMnvg86HIcw/EDhKcraYGlw6iH61+rBG9+XPxZhp8VCsY1uhm07
jTpIAYQgBGsPLD6Vxkx6DclF1zSxku3WMFGT97mWwcEYa9E3yaljrS1YFJzhD81QElk/9ekMZAdh
voB6gYv4HDbwhJlAXui5h9zaGho4wt6jeKnKlgO+B4bHny8H3zrehskgR+2K/323T66W9OEPvXci
AaLfYySRZ5NcyuhHKfHVnN0AbXL1TYneZp1rck6tGv5UzvXfK/Lax4OnWb9gI2g7s1W+XeVN7rwC
agcDyAY3Xq+Tl0F4SnFVtdlyv2vbSDzP8qeJvk8uflpaCw+B4FywwzLi1XnJvKTi8ejGPK92Izp9
VTTR++sbphvZJhbLev9szdy2UOyYbsVD19nOGpWyUVfwvnSPu+GAIULca2gJ2MVGvUdxtc7tpgji
MSfp+uMr375c94d6++PQ+pIYqkLmhOjNa9KIIePjB+EVuNmRVrcc4weIyaAEPnxgXez8HzMTDYPW
xrQVQJONZxpngUNl/vCAalGDWwJpBIGlebL5p7JcLR1RXXoWLOsbjw2ssK2IxBGP+b8ACJ2DY2lz
4zQxULGm9iarMoQ4qoHiuudNnyJ8AGPoQhBpw7uS9RbAELYXX5u5i1JjmIk1/unjEdLd7kNack1M
jZ0qMDVwMhuWH8aMMDe6cWSFyTEQqyWdW8wyB34gFMUBzu6CN6/wOIIweaQkN3zhsDNWIiNHNdN0
E8JOiPc2QhZpzctUEYFijFyoXXxBe/L8Ol+jenrhXBT+OI/RhK2vFDFERkgMiYTuptPOFe850sP5
bBeadKI7Lwh9gQtLX4lRmJAU4pmopjjzVZtV6UxelKRYFTf3fMY8xsKYv1GKRLYsYxTWeKK4RleX
Lp6A6TInjbgZKO3klRLOoDupQM3iEtgrws+P3OmlOxC1UeB3xJCr7tHZ/h4SZQQe0Oc+7gmoNGgA
SWE96k0KM6//7bP+2I5XutRMm47nMFmEs0S9d3UFaa5/0llY/0h8k4vigMwkXV28wfkEjsnZMEPO
VYvO4hI7HZ8ZoZN5AVeMiup0U6RV6nENTnzLIxzaTeC/iU4IxipThJpEH7NmgXWDsia6Ds3mK5Fm
K/f7RnhI1aI+XjbOI0vace8R8CzkkwFabwWFUIN7/6Mn2HmcQH4AdgdxUKikkJgVjBaIEalApEzd
XhmuGYnnAdnOZHU/u7YU/Mdk38MiByiB8KPeGJB7zVlrQA49abNOH+pllYSkC6BVxzh4q2eZ69pf
0K7iOJw2cginl8+1/kFKUWL9zFkTGP6TLgbWgBIPT7elXFdVOJNA2xt2TZiM/avB91anaiWqCvPA
H3SpbtlIqppRK8zKayrluQ4HR9Rt0mZZaC1z6qjKnsPlHKs6e9ApsffgceqHlpNLuIvpdZ9aJivS
oE1iDxCT+yktW4xqlEjVvnq4+64LVDTb9d+tP6b+Rg2xNBdRAXMFySaX5MTmkPd3++Edb0JKIbBx
3aqHh9sgAysRzdsvAYHvweIi3FKuahCuBhT7PngcN2eYoIPJcpUTpiq9p1OKe9w9us7rmwrl5ckH
gplrrYkAuIOjx0VJewhWDbaLBzFgAXuim7fmDNtht+t4W3jzhzlDE2Yaj0htRz4ms+nVZi4syUC1
mpwpUvFTQf39902tvBr85Oo+KraH1XmSC0axtuGCn5IoAXtFDmOMfRD8ra+qkXRSPx8PaX7k7t5X
MjqmHD/hz5KRVN/6SPS9Z+EGoy98xZ4ZY0Gjl5LnC/HHw/Wea4Cox5zg9m+bv2y5h/1oZN0Cv8Og
jj5kTOCpuJUkHdxa9bjXQ7fOnK7SvK3WZHhRWLmeNK3rAKFB82PxYZU5LaPCI5E+Mf3EoI0Ape7N
hHabgqyRXyhfjZlO17uo+8qVGy8Vk1TYthKr2glNOGg3w3sXH5RDI373Uj115Qe7Ky6kH11sRYiU
jJb4hAfNUOz+9otE2di5yKDAUDDqtTN4IuVrB0jjzw9gHkNtWWBwI93chEZWqJtr7gzzNMD14zZE
VEs9WJs0NM0EriUEXNa1d/1SetJSftGwLWLjR0HVtaQL5aJemg2VP+dxtp2zCW226mufhkkRiGTU
TERLkib+bJ02QipkWCP28ySFxumAKk8+bfmMaVcbgbj6Gd817msTw3D38RsmW5MSGJl22ATvQN0q
KmWO3quF6ZBh/0SWznoE9d+u3C0c0BaQqv2Tk+C5W/O52HH3xvQGJ/rZyf/8yVwPXxE9AEIJGYzP
ZsxzA+mTbfzij3S869TIFwqkY5wroqDx7gfnd/kbNb07eXgcIHkIHrQDMFhjhlt/1Br4/zkv/OjE
dZ0bBjWh0Biy70eJHhNSuIw5LKDbzX3Uglo2B7xuFN7D06pK7DrjqKkz3IqKeygcX+phR1NuZPk3
xB1JQNEZMacju4Ay0gCz7vfw/ol/CUgsLMvxA+R0u6xT8IvAwYhimlebN5FwofNHlnijI7cIuLg3
G4t8UKszg3hkMPQHmGdCqUHIR+skoS5/xMWhLPl5l1I69sWMJwb5fdxX5eWMGpCSeWz0ITiQ3CRA
m2HNU2DZnfJ/bPfw3aperF63qOjc9T/zlUQKElfmU4wAjsv9EAhPzkDJl9cRn2VpaYoF4viCV7jM
bxakZqJRwrzCfVu5BF62phw6f0WEL+jNPTog8DISz59Ell4iPI9sMzP1OhG4YrzZBlQmAiGoXrsE
I7i0tNY6Jk+WULBg3sQajbzhNH3XQ3RX67eBttHhIUCixYHwbaMQBf/g7p51/f0S3ZC3T3tYOdgs
7Gb7OjWAaECkdED7rLNz0jMX3iJaABS0MFK818gQSmefzbAzJXv+sI91YQ6bzFcDEfcY5+yMab1r
oVIAv8VEYiX3vBZevLqjJt21NUtsEILKFtcxBN1vtjaXpqblYyPWVAx3sgUJOx0MpT+MzR26v1ce
wX+rB/jgrJjWTvtqqtOwnUHf5jQrdNFpxGNcKCRcR9WpwcYY/ktaXGqPdofphnguOQmOLD2GafGs
q6u9elOu62VquupgcX03cYkS6hZugK90f6FHBHQtlzk4pr5omP/z71Ka4EHr8MLumK5D5HlUoulO
DNOIPUofGrDnwYNQfdtmQnPcPFCqL7h/jL/YCwRlfRJ5qZVzXgiq4E06JQw8xUl3N67JcUn/UMFA
xmZr2Kh8LQ58DtyWO5cfh2d8YOIDUwGS/m2lAAImQKu7j3cyRMcPsb0pF0TAYFnwu42+F4rJzmaO
rPv70RFrj8RiPFjA9qQF9ZAvru/JzaW4el5ERtb5Z6b6IEghD1tjjHo5rDzwptbGKUL+V0cdqIJn
qf7R3120whwGXwTY9XonegJt1HQD9BEjM29JKMz78UVtyWvrr78rvcNbGYkMrVHV1/qV+S5pC3Cy
jyqizLTILlVn7KQecwFIS0cX1oPNJ84QSSSaRxZz8VTHDg/JWkyQWnigmi1htKoK5lgNSzZc8pSx
UjaqdX9iyf6T3JXzFAf4UQPHMiROgmig0wbZVVX45tM6POa0I4Yvd1GhxkvhCuvaG0BEOOGpWm7W
K3WISx5QoYQCQrjgT4eWHJ+rqBpXYiD10Q0tDWmzD22y/UKTW82IKhYxrF0iJJ/w7F0Js55jKcIK
ja94wZ+9tJ9VYrn3dOy5FpLKkaU2xoROWxYo6i/eK1ZLa7xTeGpR0tcLCORl5expvEPxz8KHODgS
jiGDmu2YkWbRhOZ8J6QbeorNiEOjCNA5aWk3bSUEfGrAv1XX834r+LkQ/f7/cWUJ54b9EVhOCUmA
VY/CFd2z262YUG5VFJUoY8qgpx5+iDIZhT3s1EjLzR9NjpEtBOT1ULn+bhjiJvr00IqPNLU5Egqa
IAp47Arc0MHh28bidf5Kka3oyOYSagbAzQbZc9SmfxapXto2s/mkReyOVf8XpblREi8XRkkSQDXp
VVvrBZQ6QHAO1aoPk83PSD/00WvFX7O9EY4qJMvL7Yiw7NZW++ji+XLOUVXHutZ/ZNuGaca/ZdSS
kq+MMxN4la4mhpm6IY/iEmVQr1zx7uRbVcTd1uNHxB/aXfim9gFsLsDU0TkmdiFV8/EmYuSWEojC
OG7fjSQerWR99XcpmWuqpdz2zt8ddiQytukJ5LVBwBrAob6vhGzKLh9rZffKIoLzVyNnPxJ8rP0G
DzlNaHvMD+FOxl0EPnOHgmEBX+jqIWUNysQ/1fvOCpE8UT010zLvHNnnugOEZK7Y3f45s4aDRe0L
fi01q9Arz4gpI2vGd/otyhYkYJqF6+6ZzGKSl48TPSmK41U2iZT506hrlnCP6zWltU1ACOQG0kGz
0yIBX+f3Z4gqP9ujoA3+LsVxOukC75EAkh7v00zczu4/QIX0C5Yj0UxkDJ1rUKccq31Uwl6X+yi1
fAA7f/0EyqnzSZcj5MRokKu7vosQJ6hNrtBvdNxdLItRhiK0kdLofyT593rqVZQvlg6sLmdmp3SN
mrn9+dy3r76Q+M7tpnKZPR6PxVPCbfjSSTfJp1cjlnaBOFNjQJXZ0+smc6onM6whult1c0r4OZ/V
I0aBovTISwG4VaNNUV6s3ZLUI1Qb94gsmuvgjHxGLjML26Gy7RVxxU9+j83UpoT1UODSSPtnM7Sm
IGJiAWQiJt0MO1SrZvuhm39a5ExepwSCWrc8aTtWiPy083uKFWLD46vAHHu1BztZ9fKA8D/b0Tnv
TDFKkOx3141P6akLB2sZ7NvCISt1B/ERBDlDH8AgRy7zmnuetO3iHHN2xZQyg9i6Wx3KMIQxf2rh
FzfEY+onWYQZL/cprxt+O8pDs5x5y9cEnCY37/+En4YGluZY6RvWPZtBhFMpBkU5sAD9+pfr0I1X
EYgb2fmsaOUfAz7CgTk3k9z3Rf8Be9aYIfDWXbWAriCEe7l6l+Zus+H33d+Fe8zqmm/EVN1RIT+K
bkkCoPbms5EBv5spuKutQJiQvfkp/YX0kIjnnuQqh1xi+EsJZB24qyJwMPAw3D5TyMSo2mkpUMRi
y4GotnUDk9FcSV3ukrgNFFMtDO00NAQdm4uT/y0SpZ/9KUKoyfcds+Ap7iN4i865Wgo3gxG5sVXX
IKwQuZCcH756/eKPhlZhhk4GP6ZCZHGdweBnjBoa4VgEHXy/Xrfub2NdQ4E3vdCHMHson7eneTKV
kpNOQMmbpuHC8I0ffMgjemXtfHsayJKLqs2iyqfWlEiOZ7KP3pUuYqe19+fSUQF+44cjUeZjUrjf
6T3qilAiwTrvQmUUxL4n44aI5cFfvIPAy4LHb3vdGAyfzouPKUFZBHaX7WXiFhFikgvYYJZO8cTP
tRtLBnJ10V3pdL2uxqiuC8lWDcvuza533xWGZpacahC+5UGNZ8gt06sVUVbfMz14Y7mPFL7miTmv
HrwTqDsE+ZOe8ityCEGoKwwJ9sU91b3hbhFEQcnBGsa75L02K8wZMVfsJhsNS6wNd+D6ytZW4Obr
d5Nv5TTVX0URYMPO9CKckgTlNc/k9dorvlKIOA+sY2uxnjnMKGCRap+tlhewFIyKzTuhldC7mAbI
quBlEdcEzhDTm6ZPf3X74z/ZY85yxcAqlywRxK50auV0KVVsKOsiPHZE+NBUTtQWu+bDrMWKQufr
wz5+pGqsPNKZkDFNgFZ5BO7QEs7gzD2n2g28AgLt9GQOZKr50lFj7iGG6gCzPEiq23H3nKoSOxiU
VuOOoZvGWkDO6gU3mpf7GURRUzBF5ODoIm+Fgr841NMVgrEplZGSt6XYQaCeq5kAf4P9ijcHvrCY
3sz+htK3XnX4L6xoHVc9qL5Ke7WBLO1ScK3XgQAJMEzyBHiXuNoBtjosZLmuoXskHr4jaWu4ylwp
mR3E5ssw/RRuPOBdYZ1mijGVgZAAhtVj5dUEPROCtSz/32zWvJ1jMIYSsHV6p9eWJtnh9oDklqQu
QOnSIySPm9ALIltnJ2u7+yBpXeTGcFqj0WoMk3zarPvUCKtcP/yUN8FhP7TYCdhVMGy5c+AzRAtg
BMuW59KXwnbUUWfZaekXOEJMIXf0eF/AmNU3R6wepnZJwzR9kxlZVP1S1rkRj27u8GIUH/Gr74nG
xPh/tpbCoOjImRiQ1FZ5FH32RGcD63FMGxAPsEbcFPFYXR4riz+IGR6/QCj+1/wohFYNTU8yMVp5
pTlwW+puWdCgKEdjdQyOq5yncqHmFGxd2I6lSZP/O4ksbbRQEJcLXT1ULXbzB/o8pJ+TWIV9OZLF
qPiMSH4CwXXyzCVdaccTg15ivorVsDjTFH8zVZGiiUJJbU7GjpInPMON8nYJXRYvAOtiMywtrQhY
+iltv84T/HY17OU14Vkn55QbnZzdKuzUrzlm9mWRwM07VpVuaSJyEMLoaRi07bk+JyA7iSyn3CMP
CFzEB5hJtTasuCE4jfKfHriEOVySRE4W4CjRnjbTev/xujYRgPc+AMnjXBXP2SodgSDCcrqPAv2/
i7+h1CpGOimi9gST69Na//AevHqBK7rU3EZpxor3MpmC/ospGxU4nWzX1bFr9oaAYReffe/8C5Su
oxFB1oUek5yh3WLAujG1/NRZpDeaOIfpK5K4h5rkH0lAU1MrRsVWKT9lOaRvrMMONO4OOxx6Bxav
yHw4CeX3469jo6xh4XdmaYNB1rwqRrZ24rCxUW/9PUu8RJwYjsMe0uuGeLNLQlG1JZIlIf1JYHS6
BsWrqqRIt2mF2OnpIJuTheT5oEZ/U/j0VEKTqyzBRaLD87Pu4IWGo+jb6V6ojtlnZYkZV7h3k45p
9EXg4iIjsyAQzCQcjZHaIN2ES9loEbO6Z7Ii8WW5RtxxlXRa7DfC6H5an62qnFqw0tDZQvF2VD+R
j3LlOUOM0coZnN03qlPksPnBjzvyj6bPDfsjMYZEVYyMCTbRYTh1qS9QQWsUVDP7JA4ssxOjnjJA
8lP/rZKaODJjwK/OmBsel6up3V2PVgQtW5VvXeYLuI4kkiFgxVXtuofGEzaflHGNDvph3VQYTaK6
F7jba6KllsFsZyZc6CX6x1xmWdTCSv74DCxpuuXf7iiSRhXHa8ODXM8/PVsb925n5Jp7PsT6YIAK
fg2mdSrFanJViksGCk2MHisGUHj+xjJhdJgW0fKFI4rZAY9ap/Way6j9uHIaUfEHZtgVbSiBgKdr
9XuLyj4PdMVfTNRMSDnu20NvtZwU4jol0gNUpEzINc/VsvN8LQ9y9Wx+bUZ3ZVISv/dMH0D3tcv2
saG1cnDEyTKgU0uZnV41HMNUd54e8duuGNxPfjjddr48T4h63NqBqrIiEqtfgONkSE/KQ8LErCBE
o4uHdIUepa5+mh4+Ms8e1S1kaS6eux8p5RZnBFfxS6pNPid11EjcKXr5xtAbyZcRJ81S9rDQCTE/
1+7QRjeoqoNf6nXd73wS2abm9YOFwvrP3fwQ96NBBtIWtQfD+/ONrTY8l64Bxu2Cq0+RWnFY9GfS
6n3zylskDwPYA6SpL5z9KMFJ4nnQjI9ecwmv/BZA2T+vqT6u0AHrixLHaNYSppj09BBdaAXlIJeN
osUP5orWcXpDpwCpvNmZ/Fgp9fyw9+fbwkdgHqEI+XAXRHMFds8ozEexWYivLVLbCO2Tfw/Xmy3c
nx4wd52tTEz57imN8LkTNu2HTTgXqqhUzxJB3fLmuIpiFq0HReviGhNdBRC0IItVYd76Q5EDbcJK
ae0q3PtQddXGT0baZTD/k/DGKBGdMAOV6rtMi3qymQDL02/ezShGGuvill/A95UBSvjKGDT0tCir
r9RQJccaYKSHtmHpXrdJ0jN4KpjuJB8Zw6Or0VxuWoO7AW8EJMoHwBBaBuzE7kU0WmVrdzgbyp4B
OOUKeVJgy/NaTHQzdlw4Za8uxhNQ8yBPgLVFabG78Rui3dCv6R20ZIWrN8zxGFtVhXiBcvVprLez
gCKajFs6GgdvsYJe2jmM6RQYEDOSf58pdghLpdFq4bRDlJry/SKuI0JGUB91I20FrAL0+MR9LDwV
wYnJy91VfEvZd3E6WvOZsRbGnELj1M7k+EPFnJFNYOlifbet55i80oWdhKW5vkzfN/7c/Lq6rVp2
gvY2cRQkHzPb6rYwUdoyBmeg96AARUSzbGtFo3SRCO/OKvFVtMD3P0MaggkSt+oo8zR00/bHdYvw
UVRhSgwONvqFkpqMclgWgnOj2zDogaz7InzgGUDSAPoa2Xc0XxZhkAktBF/uTsrlqMdeh/uYmHE3
C0imB52Ysx5Dp7UnJmDbLjAjl+HJlVt6rTck/w6huNEL8KBAXLDE5SdOjOcAOiJZl+3hMFLQKOGH
guxn6We5+0foDdgf4r3SyooB4XKRW6t6goPTiCPjf9y+FxaXjOJ74YoV+AoQVhywE2xVMnclyrE1
6/YqRSRL8+p4UP2hPGO8FxTA9mHu0IlSwRdhT2GU9vMXYmWHO6Tg/B+1pTufcujl/ApNqA05nx5U
CQlCZSzwQERkhW5WPfcRHpjVGm+n+vU+YUXxyEYi0gLxO+rN4ZBgOvF/WFVvQPC12CEwFU4VHHGB
bH1OdoUo6WKfn1x6ig3NaJt4GXr41DZYhY/+qD2bbw7QUNMMRkP8zl765Vll2I55xCrgbOoYhKLk
IMhEMNDIv9gi05uMi8P1iAKJUJfDdvNpTnAJoOQjyeNW63cmIHhTFmB9GhVtj4Blatrddqh5ao94
9DIvSXWgF25D4f+WMdLjo4/Aj+L6PFkbVAH+Fq45jPkdzHgpVCFPSmHXUjcUNCtVfzh8A5m7+54s
V87PisEdQnfJdowfO47CsdFk5Is1nBSpgup46+UVbNs6gJ6SmqRa4S5hd8sI4yjMecmsy6TpdB36
NJYROSThpQNiJpLjWY+qAYfD7+0ehhpw2Qo3Xs4a4C1vmQ/erf2cQRP6D5FhaR5M002q4NlGUCP5
7hmsAeC6tDi3hRVDlaVsfSsqqFqPYhKjDm/dADVRTnNgg4iNA463LnDPz64+B6IT0nxDVBKW1/4b
X/wQwZeGnHvK7X9M1pa6l47UHNdDR+20GHQf7XWgYCuYLN119F0rfochSUcdmIEOFE+hIq3xG6H/
uEL57tID8yVwxejW2ylVnQ8aqFXPL0nu0mNOmMsK/1Okm8fZntzqzAlwNcwU+1lBqmJSSFUXHMhv
0RgOMBLAb8iF2DFiGyjVnWX1HBRAtWK640SAB8NT4N8zvM8ydHrleOkjvW4AkWh/uVzoeystdOD5
raEKIgXzSfxpccsQ9XGcImCh6ngDPn8kKmvgnmgc1HdCO46S18iDh59mEIBUmwUGSAamhgZi3qln
mKv4SMi65YBh2fGx576rA5p+YAheTDLMKZdg8b89Q+HqXutS7JgyIfYbrssOLweSIWm/h0UwOH8k
Ud0fjQM3EA9vcP3T59G3O2ddOSlZruKwd/yVfMOusng8eS4v4k+Bb5r84W5L/v/9M1z7f8LcOHNB
AATEy5qZ8dUgX9je0uNUKyUVvB+IxjYBd1twUhZz1kbX9O4TAgatNo/QE2Iw7qGyiW2uBJtt8/t9
kd2uE74ZdOAPRoXVXKpYakXgoW96MiZigfEbU7VlJ6hOXiJ+/dcV1evY/e6o3HgPUwNPkbP4M4Ei
v9/iu/Zn+qzhzZtRLMIF6W9fyreg8fArSuQE59xMvgMNdwlGwM5yhZ7zbOGyYRsaLIExMzoV0OLp
7Ed9oSWJ1XhCGHikDYGD99lFJ5KE++IRqr8Q88PTtS4c0tiE8iFjrRYyqJvF38F0BUfgO1o9nD6h
99CsXJTNu26iWlvmneBCLYcKI+ICPKYF+Lm4WbBOfaRPD/K5pk+LrWE50RHDz1yBWVOFYLVbVjuk
xchYRrnpA7mMXikB308LEGL7t90s/Dil8yhRUWVXFdDiCv+H+W9PTNvC6607VaC4j+bsgEhz1X8N
/zrMYKbFQxWl67a/K4T/g6NX9gzg8LhmHYuklb0r/kfZcUCV6Z5HbUX9BCNy3kHjKIEZticcpO5F
Z8dNrDb7yisLp8Gu9a8O4XM37H0zXkZwhQqDvAC/0mKXJwww4z77XJdnn56zu1ZFC4h9nmVIspqa
4YmuQvWZ2XLmaPbGJbuP08t4c7S0pJhN2CmrjHx+gaZbbDzXCgK0N9cS5s1UH9IDLysv0Xph7C1n
cwp6o4FKXNgalK5OfTHImMDmfp/X3uWQVPg0i7W3mqXZNTTNp2h35Ui8ZQFCFghAGtQxO4PHWQPD
+CTcrSSFOa98gN84rVNODaebmBAMXjgqo3impzDES7so2FJyWNkmGiNjJLT2jWylfo8qJ/b3sEdz
CK6o3xmhkzEv/gZRcnQLosC+XcNWr7hin8AoJ/eiQfOt3OtVrXvy7IE9Xy1t2Clqk8fx3Hbjz2TC
EqYOPFMKAP83m+1Ay7GU3BdMHBaCdD0M22E0gJQhhO1cBoR60OPtxDbze8fDQFdw7/FNF+UY2QHV
ZYcxGWrQnnzkR11LvlrgJaC5elO9047QgUlId4FkN8NhVll9AzhdvUi21ppb4giDbk30Tze+FKRS
Jhkp6v1UH5hqf9RCvAMlLQmAY0Jt5VqsV2hThSGutN4JNNe/X05UMq/CAAoVi5D/drhkqYTcZf6S
Q/RCfRo0mMzk4l00/T5/I1hXatsMTCoeCiPgyfqdXwNPkVrh63+jtZewKDjPM5zJuJ9HF8cwmaOk
aArxzj04aDEZVZ7U+4VqJezJBzPvPcTG0hwGPqxi6xHb5mKyig7YAkwhRcHIlPyDdfbitQmGTU5Q
xKCouVFmyDX+QA/0xx2vyM0WDAlqqQIg28ZCD6drMvm37mMNcr1XdL+ouSAl7KdAl5Ehr3rWYYcM
BRBqG5wf+eNyipHZ+MgVUQYa93uFbNpzOxW+nCNBSRpgzjSBhSdS15HRtSqZkmJtBCeUfzZUxZfl
lBx3j+Z1CLN2bPK8920uUV/rh7LKG9vMvycIcV22BftmNCZXE0Trjt/5mZV4lvj/wGxTY4IStzFW
A6bsWMMdW8trdaZeJWkDJ8kvRVQ2QBHHj8HdoLUmMQzJPuv8nzmvQXXzI8hMjGcpLKzCYEjiDSc+
GOldhaLhBqd9yuKScy048faRhulcGJkgcodE/xTN1sknSAIgk22EWToqfPAx6h2SLNZpTYOcFeey
f9j5GZUnZ9FhKBcTrjdnYLnt1lTOlKWRvpdmnr3K0dsrnAi2+Y9ZjE7XFCv5Glh1EmvPi5Ybzvhh
acx2NCMAuyHlX3lT/FW1EYmIkaRl/OIxEbnDNfZMrX/kJhWCc/qcOdbtY3UYi94R5IcJ6WYhfkaO
RRAWXo0Xs8WPWXhj3z+8NM/HFzgsYiD5N+VC+4gGDisRQbDkgII+mYj2qK/40g1SLU52wNE7+rvx
6acoHgoI9MFJq7u9sgKoBHkbPfDX8LlkH/07ydSP74O4Xkj2UXB8osMnQIAHCX5sTu+1QazICZvC
C0VxTZI+fNlgHQEGSglPAPyXrXtLoq3oJKZRM5CtsW0HqCNjGMIjHCfbwwZULIpOihEdhP5tIEpv
T1CVzflX0ZDJVZkfcPfwwFZQr6LXNojulDa1Jg9bE+wTwg9vodwX7qKrXfBEAzlFHeGVc3kjWgKs
/EG4kFQzP4CEpHUPiBAMSmjHYzivco9fK6urwALOrKu/hTv3F1JptOA1Dn9pJSgzJ5RFaHIXNvKQ
ab+Hi1KZmeTFkehVNASeNv7RUHt4ttbEiRlp3ZVq+va5F1hvrY9cQDa5IY1kz1hTCYBhN9Fwg4CV
hwDB2SBa2Y46em1j3eXJipY1ObDxnHk2FWU5SgiDXb6Ri/14zAypSjXBbnpdf1M+dmjgTat8JvJ+
aygUeLx5m1WSIj+yZ7VEZRfzxxLVzf1fofv3umwWPXo9m0V+Heq1EDs9pixCweRHsfvRF2wFWJVT
V6zGeSe/bSoL6QYQc+YpnbSkoiWgogT49Sfp4xJpnTGziF3VGQjsgfXJaiuTaMSVjWORfKQl1R6u
GWVQkQtzZ+FQis1yW3AXkVTnZDJhFEqCfIGbQNoXzrQEpVqY657LdggMsyqW0/lmyHb9ZLIEuixC
FCRAyja1WrcmKXaIxpUwVwXcqMJRmHWrUn0tLVW1PUNeM4+/7dd3VtlDHQx/DdPeJQ617kDLJfxD
uUCZGij//CfxLMdhZg1U10qYayWgLjHrEuO/LR/VeN7dK5m9YbJF/plzSeIo0JduAZWdUILL8YTd
4CFpb+CyngVgkaobF4FcAzpLgiTtBdaJ6uEKuLx3HlJ8B6XnrdBZzmSJaZxWvsjfCIUHVFXyXNhr
+JRdsFRIzF3PlXjvfLFy0im4cF1wPXQQhq0OwrA8F5R/HVU0h9fo0n16dw4cAfC5clwGSSgebWRf
Q0PhYmM3bbWUffAWWK/YIP/S58CTIufmSFjrv7ero8X4cdbw4cC7JuWEWIsa500l0SIlekBNxUBC
pkUSLsKy25ITNBop47iwEcIRxyGtlYzr+wVfegPvJ4CWmCrEwSC4WOLKbweo0adpu/22qUVDg+B3
pVkERd6mXW4Y2/wmo6bBHoG8O7/wE1XyPlvdrJT2HD6Sszb12twb2rn+TDX2tKvInTiRN7kbRK76
POh/u0/Wv8Ih6vApj/A8UTDfIB00yUfp18Xw6qy+mZ9fERtG27VdsSiRwuavbrQXPuc9PC14DtwE
ne7ZCJPhFdZmCmrVDcdHCzZQDlCDxV4B/vPN7MU9IYJtc6LtSc7GIpnnQ4bhBiWx9A0JTk4Cnugt
zY/pN//xWZu4FS7zI+ZdJRlDEAbahvS4J4S2vWYLn0Jcx8igIFH7vKdU06uWf4n9yDIbakI0u/uW
ulonceQFr4b8xD1R3gOUbzHg0sQaiJ03EiIZa0hiQfo87ufh6/kIKrEHUxJePqFaBng978bnxe48
KclgNrLv9qnVyp1XCXVFoceUTdVlZRZWpSc035L9Q/dfpODRT9bP7fFwHmhQWiYJP2y2J+8Xgp8+
NGV2AfPiLya2WtK+4A23lp4m5X2K+IEsx7oEijha7TzdJ4uzi/ytYpvKh6BSe/7OXDxqsEYQTRBH
Fsu1AGEzgSHeL63BG6kk/rJIrl+a2XYJOotbyxGXlW4rsoQ0rW5x8tmOSlmHOopr9anLCjtrvARt
2eIWfe4KM8Yousb3QXuwp6UnvzmP1FT7dd6Ow/RND4QMwy6BL0tcaqpMctz9JCi7cqBqo4PwZ6u9
KyNqVBh2+o9GEIcVWxeGz2EzcEM/M1sWxRdYDgfUMdwQFsYKqsVEHIph0x95taYumDIk7qH9LTGu
ZjmB0+omLltE371VYLKyy3CfgNsMKuT2B/2ZZ+fMz4DWVBuYUuW4gNoc7e+DnZG/vokn7aBe632A
gzw5jLo48G1pcOam5M/uPDewHECnMCVFjOXX4kkwNjRW/pfKsETjhQibDfMcLIYSvAL6/rt9RS6T
4tzwORuDgYpyIYQo29aqrmUc6AECch+Bm1zX/+AgU3XVlJRClGRQl87PauxFLK6rNAee/mApfeup
njZbFwf8v96MrT3FVOvO+pCqVRvS7A59aNDN5XUBGb/gfczvW4WiqKxlI6ibGg92j4207VniReO2
PFEZWXtO6QvFkLCBpfeXg+TQwpYIX8pzSMKgonkrqyIdOFkEH+Avej5zKH9RVapkJqs62PbkJjOY
tU78X4kR+pBMC6C02UQ56ZjA620U5aliuhgfoanzeSzu9r2hTAtAiRS4nd8ba3pcCKTh8WKOBOLr
/aYZFclBgQr2SY24poc4DP0JmuXaAlMWrD7Kuy/naBS92h84wakjzLtvX/8JdxCNYxiO5/pOvm2g
PJCMhrb/rfA6llLVbUOrYB2VT1rN1OOIHQO66nQly+rC/UEA3THzgEnnnQynt0NrDX9IHczxb5D/
JOS5satj3LLATB0nYvSWeBcnNPX51zBJn2CgUwftd6zd/cQX4Jbck9zpXphX5DhsaTvnzZwM/fch
xWUJuTJQ/NNRlHgoRlFDA7wKVbUSuvdrQ4EB9wRsgMtnk/ITp+jqKH7PXKRl8tT3rd9OH8O0HOcA
aNnkZZcq2pNpJ2D/xTF9mJtneOLibvDR3nSCu/Ur9+vtWBu/BhzVyUsFfXRBJ/KUOOR46VuVAEk9
i6blqbPXed86s5aYSi09+a/+s+gAYG/2H+kfdBfi8tfbZiNo/g2OxNtRPfqkQU0ckB6kJvUjhIpD
vIj2KvlZ3v6YXlJaRDi6VdbopCaqkx9UMBbeio729Mj8yxi9seEJmxmL5ojgRdt0BT/26stKaQoM
40VyYewA1GOP4X86lKHnAiUEiOgCJwJD7n0RgrcZHWk3XUxTJr56gY8Gv93V9S1RkU6NFmAxeCrU
ERey5ZJB+YPcx+7q3K+++S0Rygd3t97oUNIFafikwmrxxn7T4jg7bd8lgRFbt1PBrJPBP18aJDoB
sbKOGl7NU4EF+xxC9dCUKFBcHr5k2giGmP0vcorpSf4O4yAMQn4YwbXi6V2S4gAeBd1aC4JrG+bo
gBeuRepjFbBkkk1/w+eNY5lTRe6kjzmlZC+6n3nc/ULNr4RYIg8ZjRwBx41NYt45HWod9vIh+Q3A
Ex27IGfaocMsUOkSfmW+cMKuHk+XAVZ+Di0qWZZR+xO7UT1CDLzMneEy7AsEzYX5AA2yPeAuKaXT
X8meZRSL0vWsgTTBHIVEK1roZK7TQJRTEc+0c5yRu4P7R39SwfxPjntscgYt9nXkENeScaekc6rV
xkmywpHXbLQAAXmReGoTSNZihU+iWl10PQBOXZm/l5ArFPr+yFCaCW6FAuowC/e48bCwpgos6KUs
LUws0lV9jNGuCUNshEJFTBUR+S2HuNY03lXEg5IyZ97hN86kgmAA5o+Jsor6AC2FvTQ7fiAG2f9J
gXoSVTrzBYo8bYj7KLR0qK/Jh9r0JSHv/AjcjdZU7ZGEJ8sCo6JRWrlL8Obj7pxFv0RDg3udbP6I
LjNdD9+69Ol8FBVpnjsztr4AGxYs8duiCr5LHk17s5BIw/SJmUnoQKaYXJ8hQMYwVSOakqAinThv
MmSJaUofK848AnbYpyC9XWsrEZu2nfgXLLEtBbGO3DwQv+i9ZYXo4tfEx29TyCdyHcDJy1zRXaxz
DsWdplQr9kVXzdtcBgpsbvYzGWFuoi2i+gwv9FI+NwjCrrxyJWjKTAPHsnbkodlCbW7OIaMv1o3P
JIy3VN+u62WVVvWhI8ZDj1M5JyV72CWd56/MwGip/3jdJ5J9elvEaVVjuNVNItAvUMEH+c94Vk+i
+P2nbh0GkSMBQgW1qQvhdTaAIpTJvt6xyTuFvG1zAeQd8+ogRURXU/KeryeWdd5JWomu/BI4xE80
JRoHLse4dNcOETwqD9xQqlrkf1jnyPj02A0AyMU3Xws2+rAYIEIDilOKkRrLmSTk/63FKPwUCIIT
ZxisYgkIGB8WqAfpuJw+3kYB2hwYJ//cjeuFX98573C2Y/yE1spSiQQuyvpeXDrtfmLKWWbSuYN9
DsXsEaHvRvOMOJ7K3v4JPc/rW+0rJWu03EaXVbAfb2bt0zX7b69zCuVsIVymrGmesz+Qk4K0U4Qv
Q1T7ZiXTtVE00kT40rTnn1tl+0Wzla1EXfu42/n9NN/qgC4FvI1h1z96YYTS9J66+l6C++Me8sMY
9ezUQQbdtxI8UMLGyIxYojpHHc0cq5x+P4j1zRDndkWnJUQKnSNHpayZdeSbK8g5+8BjYiyGfWuz
ia7eq7buvgsyzNX4tmJYDDOlXSpG+KOf7ljYemzcu9DmSZ52m+ixtmZDYJEW8I6ziGEBeTNRAvjF
uCmrx9AwHBtXtJBrA1/3YnDOa6evaTu2HI+X+T2YlhbPX7D9ORBxZXC9i3+HC8r797xQov1EhoFt
z7ZF3yx94LEKfFJULD3teppfZKo7kRDo3Ys0DwZz/io87BnNPeV0LxKUMvto+I09b1/kWGVyv+9m
4kMjH5/CvR4wJ/zNQ9bmGDSFPSDIpAqqNBE70Tkz0t0Pr3xo3wOJRriW6Ci1bkYCiK6GVb7Aousu
E6aL67j06C/P2LEnwa+FRhfYku7PktvPCeGws3C7/ufGlMZzT7Dq1nqRXfcBdR0uU4qZfTsKxm1m
K6IzdCsYhvbDgzljRG4Ba3cTD2hn5zxvBrPZ5ea74PWbMRUHVdSFJFVWxfDPLpUmj//W87x1h1g2
JE1fi5JAaCKYmty9Xt/tj3NKfRErE17B2xJXWlmw8zoa5AMYbNRh0LXWoTH7ekWXIP2jA8mE70el
cFTYCwDN33TwQ106cpVKmPQNRLA2p3Kp6UL1pM7JH78t6MYWVevDQWwl9ytZ4NEhDiirFZW0IgyE
yv+PChpin2wr0Q7aVOZsXsiN6NF/LrN6+Kx7sHutuDUvak/rzg0SpJq7rwR2+HlzIK8vLDfhf8p8
SwKZgmf3ohE6aVA9EqkGTp3x4QL20wNSMXRBhgEgqQikSxu7TcFvTSJ6AKA4yHgj1k1oXZZCif3V
KF5Bf7BNgqp8zloave7fu/1qoXj8z6UOIpSTCELgocxSG1+im4aFjpxz2apf2O5+QBOGMZqokeks
8IFZFA+X2b5Yqc+bZA69EEevjyPyc1ME2ixIpAP7GNGcijN+TDxXIqhjF0sMrX4VQmGj+M9HWbPl
P/iGtrYx3PVLXBrnoCesWAOypCJTiO4fpzj2MJU0nWr5Hq2f1LWtQ7Vw4Ym7iuhqXYLCffG6kDhH
ZC1x2p09r4B5cQ5AdVEhVk36CNJxpGYK36/W1p0RYdi450s/okxhZZjE5aRFgF6ja9H51/S8Ktmy
omIsyuUegXJO6wcyDTM9ExEwvK269OiEUWnhP8uHAaj81BnyUvIfLVfzvpYOFQm1DJ44jkm+vi2p
joPR9tki+Aq1qYfJic+3YUWodsri+IqMSWxhWuBYG1KgO+D1rb9oLl1CjCRqcGEsbSBCdozjZl35
awIIfdFf28unFkIHBziKlihn1M3X0CTZjRJc7IBzlyq2KtRqe68WCq9P+Av7bPJLwkQSJtOcUFg1
UexIeu2ySaPgVwsHPIHiO4WO6hxbBe0dK/gH6xnxi+hZKjdy7d/tpHBt3iD1EqgTJEj3ncrt6LoB
3rBNuq+ibXciKFTc4WMAJkwmwNtPJ/Mb/SJA/NgSMHD1WgsQ6JcWAzaV1J+Z39AMphfOT/f8u1oZ
yadb8HpuzyaN/uQ5555K7gCe5l+jbUSwVdZpxlmpIck2DmH+vaXnHGN3WDDLWh5JctYlIYn3hSg4
79WdCzzzuf3MpR+D7IChsmcKhVyC5ZAnsU6K3yXhOmQUSDx49uYKo1SOPi7CmmtDyHiIt3KmYOJ6
x0xcuPTkl3nGKXD2c6GHZbtXoe7Ey9ZmDiKGuF3o/zlik3nsw3GwtIi8MXXlgwdcQn2raBwWwmmY
PWMyOp8NVh4cHA5VOi1kLumqzvm+NQ3c6qOOOqzzksEy/c76FvxsWB4tQ9Et/4lFhDkce1mnwAYP
52SeqJ5L7GwV4h9H/mAlPpC4axVcY/C9sfWzi8vKLsOApa1KPAr7WHkRlgNWGlliwaXrZ11eXEfK
kSB+5PsU9E8YsMWx8D6uZFlsKrKuAtHt4pLSPyhfQh3Ff4SlrMwoPF8RMX9JVskRvE9eHqtoui92
ZHRWL6IGKyTRuzusLDFTMuzg4dFl2dGHWjDl1ojE0ZJ+YPubkDWUppO3JHWrOHR9N31RvgFdKWKW
UGAH7x6W28POE6t6LYj3AADbXEhMhtIHnxPxQSQHJcnGTmn9GEcBHGMYQPK48zY5lKbPhcO8ya68
hOxjOm4XCLZThaHAQm5P0Fbf2ZLVppLKHjYI/ACowWWPHeZWB/bhbduqfclc8yJzpb8SviVD4ndV
Tvky2XcRsvpV9uDNRUhcH2UxJgIbAPBRNEagIZIlVStmxLEL+Le4amHLYFkYRp9h6m8pkbma+qch
8xFT3eHWrVH68F6OB3khYht7W5nkCrCuHnZzAOOfp2VZO4858vd5Vw/aCHRcQJOeBLWU46t7vk1l
ebAIL8GYPN4eAD+l66ol1K90SCyX6RZ0aEeJqNEtn23iq2ke8t8bL69dEfGBkGUqc8AAX5PNEmKt
qHhtGaX373C3damCYR5tqLk7y/D1ouEm1/l0Zz6xiinbFUZMM4kFGd1kf3snLxhiO9P9mAUbc64g
r7bdu+/Tmd+NahHo+zZWQbshFeclHgzDqbXfTlk4Onw3Y8Cbg4OgLLx8pU+x9dzRoallOZJzdTWQ
K3BPRaUJF5hIsOsv6PdwAqjZCG7wLHO4v9xMad/YMEjvY3oFbiEeYMNsh+zGodF9KxnQEyg42NYy
tJiOBqvKLydf4gQko+g09u0aFnkPWaeHrnxGtjmfBssvLDFOZqZv20yA8kUYmBv/6xcr1ooAyoIN
WWwqNwtUqlpvRL3CB3xhfr/xMflAGtp1OwCiKorKkLCSf9wpl49nQ/pvF0OLVCz0V2I25asCYwu2
3fpiCdjNU+WBQtu7e0pNLHZmkQ9vbghmoK/1HTinITABdt34jzUJtdfKiqgb/V/ErvjZEC3ut5Nc
sBmCJwH+W+R2duxH+Zv0RzNlktDaNoBltStzhu4gUou+E6KWoozxH7wLXrNT9PtWU5lfrQJ3P5Yj
I+y8u9tCbBtVh3y/HErKswVrrMKQ6GV/UsH2cPeQYaDUpGFTRv5Z9g7IKuu+tbCSzWx9WliJtgmf
BBabW2siTn8sat7Mo4fR0LMWoXBRWY4/T++VVHVzkGhQLA9kJVE26/Q4ObXnBieIsNr0ddIkAiSz
mMxBuqsnLIi2trP3K0XQ9pS25WdlM9+hAZptz98GnbergOQWs99A2NUtDcu6LbW0tHen8PNUwg0G
bFgCzz5G1UMxqcQuoGuyMVw/ss98yfVUFghGvvGJjJE01alIJL7Nn1CXQTLT6MQRlqoLU2ui+hdd
ZE+6/VD7NcZNVzCk2THPJVKk8+ECZhJBP4QjAGJZMEsOFCMi5DTSemBNObKxPwyV/QC9TH7h6cql
SqjjzlhLMPz5eRiyXvHnHCMRHe3q6n7FagcmDtB9bXqPazdMqK7imAEMPPGQrMVioCCRd1OkGJDt
WlJxj6ETE6Z6XP8PfVp3BAyLzXkER3zA5UhWr3b/bFsAc0o3nQr5qzr/X/TN1CG1wFqmZlbW1uUv
yN/2/7emb73RtixIFh/5sysVuFbNIs7Dd2kVshOXtYfhH4vQ9EImaHEtd32DhEzQ7tTSdIkv+Pu4
avv0OE9GOewVepWIxb0CGnUDdbBWkPDcb5z2T17F0vYeRG0C1QMsYpjraU6blf58Ra9GRAcml3Ir
Cd7fDK7YEPvTQjrdYjfy26F9H5N1S68EJ5oD6W5sWbYg1Yt/Ul2BOFmfAdIiAZEqhwSpemlyV2hb
HQcPS/Zqx+V/uej7bnG6p80o1iQhZ7z6/1A55GG9XgI4vri/b0zyOAZbdbj/ECqdZbgwZKxKrn/w
myLw3CkmhIGiMH5NBWp0TQc3CjgjgLZzxrtJH8a8tGIGloVJJ9Oi0iL5W90KES2V3Rgo1Pv7ufAc
venkG7dkLJ+C35QqERF5ooIkjZ23lzXxFQunsnsx7sKc7m2aj0T56IT/LyymJF5IoIznBrvQkbfd
fkP4vXucl3VHIR77LtW3cMpPQlkTaUZyw7j+6JMmhNqzWC6LdXo1eC4eSoPkGfa3UdVrdJHsPXN6
9Of4OMPlT6RbEso3JuZarT7RfDuveQlLIFrZiC721NqMZHo4Vukqf/iDlDrNVUQKiYTsl4vsKMCi
bl+uYBZrDn05g3nkzVi9SEfvkj42eqa5S94Y1W/9t/mdCJjqiPhrp8PtjoTx6kLiMDE341LNgbnc
pDvUhdF9YccXyNFArVqt/QozJqm/knhDS4zNpG2lSpWjSe3uktg9v0gafGgqNcGWunhfF2p9JMfP
ZmuY4TsA8mEGVm+ooBCMxbnOdfzgLP8NWJo8Klwn7ov6Qvutgf6FJzCGZYqXnItFM4PnPYoSw3Q2
gEIqcsTcjKVwYj5xUuousJL2l5ZKOYVZ183Yy5qSWCLXugMIPMFKeIWoT/caK+wuH9kbizKAuB+W
NaKz25EGfcUxOcXD3oCza3s24Xhs9XRkd3300fYvDo5jf3Vby7jDNVeeGkB7722/+H4uGaKwHv/8
Jd2NgoErguTv4j/S5BpjXFn7tgq3ZZY+Gnrvi9S8JXKRaf+zXr8iT/rQ0ObrL5SI1YBj9uxcfkpJ
cEKhiKMgYs/pzT2lBGw3ckfGosNIBmmoGKXUQlhQsOkJ26iPNBKPQge4h5dq4sZRspHNFdX+oH2A
E+M23khlQnxzO/f7kmJSCCz4iT5IDKVkPP//eBBIvPkzVGR3xNUjKRP14x88WtYag7t+E6YmuoK2
kEi0A+Emi29a9m/Q6zc8Zb2xsiWdjU+X16LYWldV+sgFxNS5y/+cIdsze/0Wt+U98IELmYtNPKdi
3y3dPSTLClnQlOIDXjnRTRqRyE1lvXLkIjwm2jUNZWwwn6BVq5Z7iAdpq04D+1Xgu0tCWQqA2/5v
QBRLWmc6cOefpRjmh1Q2FvfFLboHh2RhCLqjUyXJPBYZfNGk92RHgn4vdGlPU+NSSPKgUwwGytxT
38tXP7pIamuZthw1/c09LjoDjAsa3fkir4gY/AWdXB7Nnwhv2ZjHGwk3NDqGH3uTuWIQHiBjFwLK
Ij2SgYspZ9WUnK2OC9VsQcIuZ8cS6wS3U9VaPcxgBOllt9IrzQsP2u3CIVgz1zFJgEYbwyCCKSNv
/SrpVnxqbGZoCGHgDiFkZxvakXhOtWfyfxhsmydJSO9pCq5HlHRV8o9mGMMjq9rUvZBP8jjgYQ3r
mGLvQJQe7GXD4WQjmFrWDxxQqZaOeBHI0x9eOHiywz5mfge3DlryfkyZAdhjsYPlOhgqxLseFwZT
giNv3305CuNWInkQOrTjlO8m27+w/x/gw3h7L5J/bqfzV4cfg3hUwFa08N83kI147TwqFzvOJpMY
XFQOb10I7OLT1ddudx/RKwb5LXUzWrrog5i7BcVMMimZ8eH2VGMCUbbmWjpRx5S/05R0/LlLgyH/
f965edkPDE4HNzppM9f7w3CafcAKuO5e9fw+x1bQaRpX3Slh9ZPPCymQZtgRVMpfmXy4Svw2XJKd
LcuYyS6Utylyv1PLKAJC5tJA6X+kH4JB+LzICvd56DTUahFp72DwdxApAdJdOeOyzzAxHzVf9Yw6
okCWMZvy/YCPTA27s6no6EZFTZtr4qlNXLKIf85HooMc/Y8rnAI9QQXpzTfVx8qpcDwzBQBFXGFX
smcJqdoQt7QqOHpgAlNXAGs7XEHmrOFf6W2a7ygRULt8/WoiabR8XxzCpW0hOoq0MW8YvOYiYa8p
ac2NnmFwNI0HRohFbnbnD99566/39I7tHASseZpNdQdSyK7LY78BHXyJ+MWRZRl4whTzczdYz9dv
3iG+A/r11j6T4FqTGg4/gOYREEwwbsIztLeMqyxO9qhdFRq1kiZeaafLYOTBSgo2osPdljOhMZd4
LRZIt+ZjDnhy8bMMVguXvnDvI/dXFwM6mS3S3nPBhw5+23v2ADSGj8+0G28VkMbO1BpWSaI8q8do
+n7BwbZojN294UZ+56sIiPMVLcsK2RLncLcZCTJ2GMyJgdv7EFhn2yLfGooDOE8U/7SoBC8l4msZ
D7kgGPZlDJueybld2Pc8nEP6AxYhtiOcxyWAP1Q6Du3lfaklZLbXKkt2EpB+I8hFREVCfhSidRTS
aLGzhzOzV1cn9c3Oe9hX+Bgl3/bDcIxkEyfGKztwDBu0Ko20E9h+cXJAJMlIqWmQJ3kc4D99D+qm
PORa//Z6woVF5cSLg7ipi9OVW6xIVLXCEXOfrPWKmIleb0uB94Vcr/AYVR4yj++yTmVg/ZdxQLvU
i+sTBHxmOTRZqOkjrndeNWUMG1JU2XEYdUBCu+sAcpyI4MiQPOT9m162zoAl0GyGNzBCXlLlS2Rz
pr018QaDki7yDOwotF6u3CzY2GqVHAafOrJ2VcGt8G+L8MA5JC2kZprsiNqHUbsuaOen6isaplpH
pdpYSVelHkNKEFLRZZFwqQBvkDR/t+/nbnbBqoBAAw/rfNSS2Yg/7jtikMCdyO0kvj9DNrfw9EIq
LZK6mBm3KTVbY74s/AglnrRVhsOuVonElSha38P7lqjTJ5CrcakRjpRmM3uMgOAhvXTcTX9k+Nkv
yq0O2Zq4hVruzOd6+gI3Xa/sfhUvyCMVq4UeSOe9XPm4yIbiBP6huf5ncW++TvMmfiIvCegGL08R
Vf2pi+27/N4oKyl74KzXlrQIBhi++bwZUq3HeI7AQ8rOTgTtc45bV8StkYch4dYk/qjRh9x/wkNZ
F2/D2rovuRV8czSXy9kEUB8qC6NkPnXWduAljHXayERjvUw0COvPNFWvNCApKrqQdZmD9F6O6NwB
0Wk3jZKlRchTowBFmVVJDJ0IdO8md46YAOYBCGl5/1bpTNUt7RxBLjErzDG16qvDXSQi/nmpC/59
iWbZ3wGGDh/TIOgFnCL6SQKqb4D3mMQ4Qt7wbA5Fm/yQ0cSvFu3zjjpiVqaGGKhvCH4nB95HFrXB
llDyg74rT5f3RBlwxDho6Ejfhf2kBIrhnPEQLbkWU7JYSp8CFewSWoKOLiHVt5CsatJJj99kSebc
bu4V8BieosKm0EH/bjN2ROitoPVm8uz3Gw8HV0y4I9/IlGv8k/gxjOK7RX4twjmd9sJt3rCD2P1O
l56qMtam23nu6p2A5daT8KU0GXtF73nunQ1rTIxzJmuH8KlkIEE9TYxiwa/NDeJFoxtfwRS2QPG0
vicQCcOE7rx0tgac6CCXyFw9f8lvLnMSQg7slmX5Kg9TiiFodtOLApCes4ngyE3YfNJVmveJx3JT
bjlrx99ZspecmAuus/Gaz36D+kTr2BokuHZor8BAzKAnbJoh3mSD5zFExGr68lsE0VbXXSwqAqZi
Qj6E95kF3WFl7RwJ+IlPOZCrW1l9ZyI+H7TwqEVQl3qIvC0oJvpAKBRGwQGRbFrSJJNrcXXtks2o
MNEvpxG2r2/mSPpGFNTAluQRtc5dqKZwfujoJwc3yvaWW7Hy+tHcSTYJZJwoU/y3agLIqT+qh+0Z
rfP3TWj4KG/k2Ide5NxcB/2ILaedWmf+jEuPkrQXpIgi6Y0ie+xApFgU19WNFmqWQNlXih1fjluv
+IpKykO1yEzY1EBtWFt0QfgNm17yqcDLaJSOePW7mODXCXtLZIGn0DTmqvyqNKIHPnBft8rJd/6w
cpXc1fd8XV1Om2Jal9LwkjNa+IIH9FG+l35y3nU1ZKBWQYjifuig03VuHR26tVu3YTJhLJecX8/p
uOeARP0qP3hAJRT3VgMsVPlBRs9n5jionZRDVxjvlfbj39OFojlsOTrIEf6g0pJYgmOoLUBG4Dnn
ZqytzCY8mWcpSnI1aGG/njyi1eFJEvrqk+WkIfq+ozx5//ihc6zHs9TETNi+d13/keXEYWJ+rugz
qhs+00oS+o2upXVz7oHdBsg2vte0k2iyAH04SrkUk/eqvwThVPEa0feRTje5V6uWwVv3FfGSCjYt
15dwGsPl0x5iDNbDGaRTi07w3+DPlNXRpremckAtVKVX3RkObaBRV981uIUSLWmpQRo1UL0+Gw7f
1eHaQepSXaRb7+oaytdHneu3KEuX+hXTAOZpSIaLceQalzPWTuknDyUCP/lhCId1GHduWM1wZYlU
IAB1r/gZgZiGUMAASatE3bTWxxuVnjjFbwdY4twPq3Ef/KgkAjG3qB8t4eP9emm0TpUarH+lpUuc
rr5CYEyIA6IevRdu3p3fKRFiRAqWA9n/EhITjSGryEOOzLvQ266RLhLrz89Zn5kTqP52xJqQt7Jy
aAnmfH6J+ImS3j69e1HPIzoctIhF5K5sMBKCDsDw6xqlS1p9yJZhjwGXAhu6bvpYSK9EwOdJbm03
xX0kevHqPPm1tDyxpgFe0/zuyDrCKpLKSF/APnB38FTnvWABnWTNEVRWzploPH7m/fTC3jEjxqOj
Ddp8wNIPpzRNeJlo7rw/zh9/gyGPvW/SJJaBRFrbZsBDS9JbmDh3P5P3N1ELW5r8TPg5wruk06vS
OJHjBxSqkDCsQtDV6xzW+rKfBzvsYxLRyHcUFxz+ah0fHdUKrc5T+BQyZgo5eIla2ccLa9LCj3Us
dUYm+XJJG/XP8yHu/KKW9PDEnVnHW+PMLPE6vBDmMMS+CkREyFzRmVjSSRUk8rrmias6875UIZG7
fc4S7jE3/w7zNbz2jBfZDpSbRbzmJ+aHJsTHdT/k/lThT/g/UmIIb6GBkyHU1XYMM+N4VRsP/KJd
GkqsHWdzZzZPtrVqEealSIAv4mXH0U5Xk9YfZ1zkvYRqP6oCcfwsVovfoUVl+dHQ6Ij7T1KdI761
n0b0U4iI33t3UVSIGIhIX7WMdj07kfPgu0idPBXPxtj0ky91w96EQGv9lFLNWbQFpXxstbw486d2
MYM4HgafwhIq8bZFSrf+5RCXtoZPv2HcV5YW3l46Ma2QMilC9YaMBxr2kkbAkmZkPcj1JC5j2y+d
le4umyxEkx7Huoa/iwH3zWybo2bDHOa4U/+3BB9a9gsN0Y1iPq6lw160Zi9tjpo2CCRkI3hBL256
9iijYk/0gvOgUt5kiI/Qc1YvJKN2SHFHGJ8dpH3kRX2ZRuYlAunxT1EpZbvefZFI9UfJCDXDMcB4
42K5bkEYTUAbJqc+cVi6UUItTJR+Pv4bWAeHHI0hmFkt+y9GRHgH9U7Fwiha6hXFR6sbztpI86tn
ZKM4wmOqQCEebRWgl1+j3+1nPqKHXm35s6PyN8uJh8wcyRSVcWgtSZlE0T93T5VKXRdYBvkC/RmG
GF4O5/7NFuT1ntvITMz0I7tPhnHEkjaLJ95pDXKJXNemKnLw2sZmHNq2PbOIzwHDK/bGbMU4xThP
FRPw3FXRU7INcR60Z6/El29Qa93trRBC4yUZ9dfgJsM3D8pieZMOinBUAIMgIb9jA0t+UuyR+X/x
+J+BQitL0v8a8aUlOZLY58BfsXrCN8P7Lq6kDay5183lMwbzMzj44fkQe0KDy90aebGxaqqfFUnx
o3mOsVQIqiU1DiWbAaI3BlG+k4uejpIwn5LBni2vvNFpSIF2VwgiuZ7FWgEZ69kTXigCcOQKe+iU
vTLcOHzdyoa1Y6OxLBHNNydkF8CjOZoYQuA+gPxVBNNr/82FkGaddp6KVYnUJY2cMA7po/s0kztx
LI0LiE0n3OqjUYDhKbuQig24mDmT0abxAl0wyRTHNjSXIpfAm7ZZSCHUnC3s320Y+GjbL00vE8A/
aMCW9ligmQBA2Xfp8+Er+nQ4p7uj4DiBazeJHoaR/stlPvIQ40Yc257xSX4Kk8iolz1vqbwjclh9
bWh06CSBufSGWPLvb20eZuNshptulUXxGSNenPiaGRZrXccRFZTgl8q8U51V2KJtCa4cKv1ua/eQ
Eavh2aXTfYB5Qfb3+bo3qehyZyqbQbHtKzydYalwKZYpvg6QP/YgwtgzvpSSEKd9QFvx2Hx4y1Ll
enWBwxGQgbHPUUxu0eO8LI3Co1fz0JNh+EQDZhFOjKpa2oG3X7XIMKz1rNgMTKmtbxtfuc1fOILe
Uxd7p8UmiQpTD92Mp22i8wslfeLVEBP3bG0a3OXNIeL7n2SZVORGaB5aWcP160LJIEUditOIZdiS
7itewdw9DPjM8D3n5p18OioEv4hvdq3kPRYlsS5dR51ZjjoiNxbuu+hc7bDQ4asfl3zl4v3PiD2f
H57ytndEpyLixy0V8Q32xUCcEU3HJYojJkzJ9wN4Ja6RX3SVHq6AqMnUjXQEn8CTd275873r40xO
DwVBIWQk5W8ck7YR45kV7uO/8ATQ3kwgm4dm08CV+6/sN6cXhKgm4/e/QQUdLu1YfjRD/ENrEzi0
uVafVPA4zBcelYLKA1MduPoaUvl2I9F/WNqoSqwrEP8p4p2xR7xy2b6h74AjH4SCFnBtzKVKptUr
xirjBi3xe3cBUHNGNPb4C/fbFf4CCU/FMoF9nYiOOLvT5nTWBKsjJ+hfmmctsw8oDu4jyKOKwQin
Kk0SALRJN1W3bNjrij2CJuHRHNflsR6qQIKgI5P8/SNr1nJlkRAF9SkBkmPopMHIANAIsJxTo7jr
oNeDaCJJlD9CYNjdDLIZ0LLCBcmvGsFL2WnDvCXAEwxxv0xTgDp2lCGLoDDpIt7iMNgaynH7lLkQ
p6iP3VyGRyurKVOC6Kl+ytDg4p7NuF9mtWHHPknW6Kccctr3jZt3iuZAhdxrt6BwLGD5aBCvJGm5
Sq7VGUFI5OWnSSrKu221SCwUbpTOrlGtGHGojpAQ+TY/mQpXRHCaYWVYGdyXI5raCqEq/sjcQ8vF
zTsf6T6ohKepzXckTVB9wqx5rkvvDTijdE93Yga62E4cApCvlqhzk3AZ3uE2kvTZqdUb3+MMQS6r
ETB4beBcr+X9//z8JaEJlwRZXHoAKE6ArYEExT2axeEolwgdMsZJz0RaMjtMxsaAuK4wLLeSxjC/
UCWZbj2LGnZGonH+mBPQRLy4fD3NpFaLTuZ3bD81Q01K948glrlOjosKOdGVFkNQcWSegMm20Nx4
PNipcBVIfkblWwGB+J1vW2mAzm6lYS9cgpQCoamRkY7wm3NLe3jpNZ+yz3AstNcT22sjMo48PTKL
iNTIthNDraat8MLdjPF937WJ27EPw5yFiv4/84uoUY0/OcGhwa1jXJVHf6wO9lG6K+0LFg4HttZp
s3JkklX/PJVUNYMMmKPjDzypIXKicVyuv3Jk+UIj7sW35oTyCXTlugDCVdD5+B2ar6YU+D4Ooy1B
U8XxXTrguJ7LBm2xszmybdFqqsDChleGFYZfxkGng0iZEyxpNZWQTJh4Bpw4bXSypkahbM53xt4y
/G82AxZJk/RP1bBrS89JMeXBBlj2oJeIpFO0Xh2rsQGAn5cEbcs0QcQVIT+yP+8j2Fly6ilq1e46
nprwu1NHFzxl6VM+gjKQxs2BphqP6ylscABr26JV5M/8ebROinWXbOmwCl5Ob38ol8H6KkcvmKUo
DRVs/4tTcjqY9dUMneN5qkXgc1HP9e1xHSHE6P4dnjpx1rMst9/BpqjdAxhS+2wC7ntRa0Q2H1zp
fenO3eodoNjS5vJdRPkqMeo5caFjARBVERilEpByUW/YLjkHUI2q6e4DWb4e2RQiqfWqSyvwDk0x
HaYk0DaDEyCyRinMXWMXbeTg7GX+Ec0Gj34Y5D1mgaKfzCy4P/4BVBqcAWAa8Ik3vWhqV6Gs7w3O
s+Jx5BVZ9npqi+ikshAjNy3ly+um0JuZKUzM3kAgsOCYsArCq/bZzhAg4nb+oGU3KN5JGqhikSDd
ra2CQNCeQ4prVM6mgUoUre6wqY21omIncumFZYCtkAXVxCeVwTu/uY0+Jw6H1TQUjoHnf/OesUyq
Quwyz2mRPKl7YeLjHnlWS+7JvllfUSid5sFhnfnqhoTA98adlBohkmLWUzlvKIN2VZLlh4XHQq40
z00SgavMFpFHy7Nqu00Nz2piO8h8C4we069Y6t4yk6qka+1HfrUOvXReKs31lDRsIvcWyTDKuZ4l
P+pVgHDW5yTQl1Itxm6ymv89HI7vD8X1XbuUTqMjVW6L3tb8WlGnAiJHNhHILswYTAmRWAYyuaWq
RofoN5pXUSPegR1tHnO6YPkLTgCG8vh8NHqU3D/Gquf70LAQcSL6T9tRdc6wppH4YwUxymoqhX8a
eVZxg+toDyxePuKxxW/I4zeP/IuJj72xz8MnKCtfNabrHfr0yH+GzzcwDBRyjm2zVHT6YxNRl8Zv
pgETe4KT2X7NY0RwIb3mvAGv/Ro9ddoNWZ5cvLHQ4O+EEf3/duAtnYqTWq0Aw66yFVassvwTL5DG
9NCH2Tj+HdlC/LfEt+NIoZP7Fv1yaIFkE6ZJNyg5YoFWJm2KCe/uoPQDrLyExKtFiLnym+sm+rBm
KcxgJahOPkNzcgkcVH5Um2l9Bx8NggP+qApNUI9RxWVSfWeHuQkL0f2b1GJIZRNU+GrqQsfIkNdC
u83dA2KgbNGmd9OMIGsKioyAM1MhY2ngVp8o5GQABQCnKmWTgNhgVComysLl4QwJRjeey2gYMGX/
3/utVh552XY+wSvNSoKoMLRe3jBUrK2/vtM4hXA71HFKrxXiJ13KZr5LUSB5kZ7VNbAxvu31Nf9N
iG1BuSs2lr7/8QvwgTK0Kac6zf/wIkMnW0XYKMNFGIC0TJVR4PNKaSmEpLiQ4RQQIBQ2ItQKLDpI
nc/ygNEAf/prRITD+2EbOQyFzYN3+5mElVS8tG4z3LxZrtB1mIufME8ykWvl1yLfwiVI1cJZX4No
qTzAAPP0yzFTEijhqBjw5QEBwlbXwG/eqeSTcRxJ93YUV31XBsrk8+0ETl+KpumrKoUhh3ZJhIvd
opqqwyg9CEg9/kadw9QGz1gFeI8DvfYhPjCu/2WwxYWtddYlEwqVjgZEQpbtlJ56yRY3Qd/BrlXH
qxvbh1NAXxkDlCC7IdDcucy2l5OAIHjpPAakOtuBiF9vHm4aOProT6ya2Hf7qTKHfnkJE4Gwkuwv
f3cWCkYtgeEDu5z2cWRc3a0ke+hFdd5KDhVt86KYzGQFQJwXBLKzJbzCXQqqBvyqdWbE48LMRUz/
qyonrK0b7EP5DxCPZzXmQo6r2DWQ/d5E9WTNWYcsqca9mZfmUZDZDLyeBHdpoHbVF8DRvR0UZpmp
ekfRYjw1CCuL9zOedG4LM74hZnUg5dB2aDTEL6q5CJwZ/WKx7l2Im0pTb4nR9NnVohyw7NEcJSMd
QtX1T7xVh/y/OEeFMUmI0WwLPas7XubDXrE6NZbmN72pCGtBLKCnQOPtbZ2gzugnDUxZ9cTV7bQ8
lNr1a/RwwiR9wKPPNVwm6yHyuJJ5GKeHAQdSvtyO1tN8s4OSdDGExvQ6ophpbY0IfUhJW/ibl1Fj
o4kxcFFYadHXJe9329w1qi+HJiUpPhpNQown7ocNiplHBKfCUTGvB1rg0xZGn2bfGMuHKfO5GgO8
E9MISTi3gEVNxjHT5pfllt73KYp87en/2c6U/XW1aC6v+46dk4C9qnHKKiCVeceGLLLpm/nhFayU
/4Zhv8s9FAEfweBGDiLLsVwuF95gHa+0XW8z7YGDPB65elWeLekBQKPT7LMCQjWTicDl0uOMTIcP
gXue1HYfGjPg687YnlyQg4kNdxXFUB429nU91HaPpYNOsQA6o2EibMm6RTC6xbNqA4CHUFIdZPtr
pcapBpgPMkRVxvuSMwBzuFqPYcG85tyN72X3F7kcjNaSeYINpBYcscaIAUq/b/3Vnxuyp/9vrBpb
Wmrh+duS9CcjpGB9du2RfGah1DuygjNOFosE47Q2hr9QIGooRGW8LpDGptcuhioAsme13wub2vAG
v1MrzVgLNrZ0fafk0qR6HemTR3473V/02LQSg6f1PDS5+E7eWXZVBp9FJG97HguzMY5kro8Ksl4+
4AIvbrZxaI7U0egOe6/6oDOLj3TuYwHc4fC/IT1pQFliHcr1uTpn7KXWLTqhcApx34g0EgRBxz2P
81XZgxPzttIQCC5eXRtLFOZXkdiiKKEuhb90ZsUNFXtUTM1EFigQ5zs93uMrdw+WAZYyBYjdD9yD
6M5Hn4EQifhqmd4W97m6l/92zIuJuRWs7qOtC72EpUPTO34VbUYbmpPqm5IXyXgA7vNVJERguu1Z
Z2ZT2A005fDs86SujCI4s14cP8JtKff5QrivxPCrhuXlSyJ0a3amWDUzrm7+fuVAgCOh0nUzLwK4
UVgNUAq2ycE+1tDt6qDIbNcOJRl32AUizvkrIEgvyoHlgSKfUYUgdMgp4AKPq3CkLwkRtjlFDmDe
ul2bpKEjQzgEb79MReWFGdlvwICOLUnrZP+b+FqqQOgClsqcl0qRau+3n4GPZfyS/hxKb6tZpBSa
IHbqRant+UKda1/4z7fM+1DeaCUakavxil/VDHRNIoFxInGKlL/6kv4eiwtWHb2jFpLUX6X1GtXm
0YuvlI1MZ/Kzu/xR6+ujyncuhpTay/ogQ4vWCt5xMp3zt4ZPK2o4MiH8Sw5+SUaHBX0xNdmx4beS
WeCWlANg16NTMDuFZkfdt88aSYwpc2x7EzcesVw89mWnhrJwwP80tk0S+WLXZbcQ9kWq5/KNOOG1
IQ/V/u3vL+yHTAEBPAZBzK9QcdJxDnPtZKiDu0KZr2l1J+e6L70KFVd9pmOiKdwceXG3p62dK2Jx
WINcmtmo7KoVvYSqB+3zQ9zWvlA6ffoIaXUSe8rL/hveQ4hzaVWHsum6WIsMlNwQHoFI8oP54/w0
kUIYOfBkMv+F2vE3Z9PR6EhPFcIWtki86tEh9N6k6pMW3fbuzDvaL1fUDxVZt8obpoOj1an1FpkE
Lpc1LHJsoff5MLrQR4KYCO4we96gl4RPnyi4dZb4vNJpfl1yMIa1atjsGbpblQqLtLYyqeww8fUv
DlYl6SzPp6bNrwWgxuYrRYOuxWA9u/RW9MOQ1Uudoe63ltVOFAq0UKJLLMRKH/AdJy/lrkzvV/YS
rr/elo3Og64/TdK3/lWCchBkB4lyAeUi51mnexV0IMr3/SXC3EsWoyelgliKR9a4eAsl+sZ/tynU
mhpVa1oEHNJDrYFBoCjxemxb3IgcNK8mnS+0I9LmoBxrTAe29VTOlgfCrELmsRKR9nmSmBoy36Ff
AbDhPO8Xs1Lw7YA6kKoLqet8OREtNlp0Ey1CfqGQCZZkH4d7hV1T6Yuu2SBcGa1RTbwbmKfImyaQ
f2lMtYy//OhucgfiIBTUSDTobj4rXXK/kQktHPDXShk/arga5ErgsuCA0IMHriNLTFNgFh4rzLYl
Z0tI/WM9rM9DVC6BjXon3rw1lXhh1KVHHIZwvPVbjLb6cPXQ+KotkdDFK4qsCfMn4ScnDASqRb9s
WdEVtE+vZACl//Qc/FT6jE07swIiniArO7ufnO+GBRhV/CySrsy/SUPWEtcJBjfPAojp/P2tZ947
KQfixADqrMnnoy3S6GM5eyqr1uZXfsWWFcstZc53DxYgJp4ck1BrYx1qejwvKzeoC/yx/O0w92Qy
EcHHOJF1kp/YsJkN0eyvOikQkwlTLZOl6GtZmj2gkebmhHZ1wDK69mzTIamZ7I9ARuPl5UhGf3qA
bizXmnVN9reABZ2KtTMuGOBAH9MU9h17ZOlxqDrZKEM1fIK/t4gQiHv93imTbgd8yeylGaVtngji
WabJWTUG/7s/7Cs79i/qd3YQRdisn6TMy2MRJIFjNm2oBf0TfaW1+D1L2fTJY6G7Fv8XgzB+QeeA
4J/hUkvzwybM4dYgUXSkuVowF4UTprKcWstfNqiD6vEhMt3di4l7fpvVXgX7xIGz6XUUUom5zaR+
JU3rUiiTVL24nqyA/jBC2IVBUNqAgl7dNsyBxDVuhpHNSD3msAPlWm5UaSYpaji1PizUZw0anwOg
SSwBGDmk2/a40+pRodl6JLbqajT8VEFy5fuHtLgiu4jrA+IK/HNiTwi3PIDH+xJn+/aycf4EvabZ
2OiYygD6pHmjHQYNcT8mlr1AaNYb4a6re/KRGa6rAyuc6RXXxMMQWN0K97OkllFEiOibY+quVh7A
rLqVtNmw3XZB8ZhX39y8ah8sBUa4WsD6VZHHf6UqBv7PMwUrkEzVBWIygKzcrMeBWy4NYjdP8S6/
b9D052ABUKaIqCnL2ruFqndjlAUR2u9fipptICUJi6UHDfYVLdOTUnjv8IPkdxHVUKSu0TB1LFuf
88Nk/amrFGP9yCq04ZdXCUfxI9c8LpQGg4PXX/wKK6Nuf73tL8SSvHHJaPPkcSk3c4iqcP4wBqSk
o554A6cOFhYL/GYKikUjcG9PVArBre2Y1T6yKM6UyUmvi3VrH/3BGT8pBF8NKEAdMV61hsnQaaVt
ON+LK7YPp59P68iGzWQ7olKaMiCO3dGZvU6SsuX69GyqEc7eRDxxZTfCLU6Tf5oEP3iOdfLggevF
tl7+iHU/0+ATi4Wt+klGpz+D+zA1Qg0PRIqWgh+cGvXPBcdQuueSx+9JCUSDe93hUHRclF475BcJ
6+Ok+g9yA6pRzAhJPp3gZgo/dJqsuwGbQUyP63fovgXrZ5PLHgArJJHIX66JQB4x8aKMrESemeVG
0lWhlv6lRtqnu4izCNkxNN/f93Z7/+BB1/ehWtBpPi1JE2agEsyrvv3P1cZL9rXffCmdLlLGqOe+
loxe31uKFcWJafFwAjpAonPVuzkkKMTLYjbJT9iEiUSRwJ/QUgyqGjTUAbaB3G9DNVn6cUnLguNM
P9E2bgzqFL1v7qpPeHK3e+qbCyvlKL3OXYlVRijw/39/e9k8qK6TkOzVbA45Zx0480msS0QIEieY
NEfT6ERSgHHO8V0YOsramgZV28mytIEx07q54aHS12RtCPaUaS1094KrffRTTOCnMOxR4ObDiBZh
6KAC88Yp1vwH85hF9uQkxfHP9x1L0J6BKqqH8NGb39QCteAY5C0dQ/D/f+G2XO42Aa1VrT7G5Y5z
rebBHbAWSps9ueiteAnSOP3vedx1GedA6b/ZtVSMTZ7JGUkBhFE54rH0Ga2nh6abIi5rGMvLmnkC
I7RqxmtTJAnii/q3d0WeBoNDAwE5VMpF6ZLEQ0+d8zIAfpA6V2enVm16ncPVj0SnXwmcVDCmRafX
ql6d2tUXku13OoljsueDQH0iMSSuys5IjzkS9S9s40ZrG/sLm7PVIAvW2ACZZbOORSR+djDrC53t
nyy+l99760tJODqtMfGvd992c/OgZYc2EhsWYET95nARb/JjIdkKUdiBrBp57XpfhkqPj+Pr+t+u
tWzLqC4RNSGJKew6mep79ehw2eLYUln6mu+oIBSofQZQFxVZn7VhPNyPcIlmQQ7L/a7im962Pryn
SGNaLE4pj09i4FMird3kuhPZniVDBW9QdDN2IFIzIVoRUcNgs7QXuBQo7qtdwKmKJGGHydkNO6Wf
N8GmBOGBX5SlBA7R+lr7dW61CrjsIQKDJmAyqxul4huH5WcZOogT3uWo4Cks2kRSbHLjKjO6pebp
XAAw9L0ckTtXRA17yaOlWpQiIe9vhUlIsYW+7WV9oZ3LcLFoKRuqAVieuv2WO1wHhHPZV7i7+xgN
YxAIczFjDrz5IluEkfCqiThQ5RSIWyPYcplP9z2DKBfqcDq4nbBYzrWDvg/pva+lDmQ/EUI9mjbJ
Ce5ccqfU8pQ8QbVFbG8naEW4rXITc/Tw6bCF3BUwq/3BK/Y+bHkJ7EXS4M1dY+OTGmlP5dnHBMHa
wQVUc3ZHQrrxgGm+kXfE1XJtboGjcnbTExOQ6tLfHlh5HvDa4h8XHeEaECwQXZxeFkXgwcKc9yoX
EJtQW3dr39aki5jj27Bsx2Y7hRWN8SodQ5yJ9CzQlobSHLFMgYsa6j05PbksWK1XGH8RPadBNEjV
+xhXAabtjK8jn8uJvytwcD2D31ztwVKFiOHv1cLnTjt8KAqyiYRACke4G0YTp6JrssUWNtjRWSMo
0duq467//Gywcg/Ptb2oMatcWOCBDYVC+VmhcM/TBi4oSCIQRhdGcedfqO6YTf5zOPTPOrqucTBU
lJrTlbplCq/V8lk/AKFOzk8NbNQo1kiGsmuQ7AW3ztTQaj4G+PBUpQ17Dl+JAZqGjnE//V/1fK6e
ePPvuOowhil1tbsUyldKiRXkw6Emrpc6PpK/WY9dcAE98HlKqmKlcH6ICMBkHSLVRMPtvM1xwGeu
y7x4ms5Mwcow+xjwYKH8QbOyIHAkUqpZSJ6Gh+SIWWLbIM9X73lCEM9FrXQUVVsFkLRGQSC1YfLP
4DSzuZr7yGboWv2Ytu9UqPIEqxBZlmQ8g0vbskNexJlK5cpf0PkBpet2+vuvRPunZ2Ds/o2KMnsH
fUDyh2pv7nYZDQm38TYUq5Nq1BMiLuqNuLb81jjsCwJbfrr1EdZLjdB3dcABobCV8T5/EAPYN+/h
bOFWkNzW66h8ItDOdsgIuY6f4SCtZC0/fbFl8PkA/fbHdWwq6mtzp40xdiIfEQm4GFvsMNiDHJVb
k2zjRK7CF6Xq4kEiQQ/CE/fSDrOAWfWhm7uFIx1G8swIOrHSGxCNtpqOPEkJw0gVnzFHK/tN9zO7
Y61G/9o4XHzQz0A9OOZDH0qZUAmGKYGE71Sk0+I0uKwdM6xY5yJ3Fb4OWCqdvh0n2HjH2eNQH+o7
BNTrbgxVfbSGso5Gg/qVKJboiCd3D0PJtlrL48NSdcd0tVyJHlZcYu4k0PKk0PiEcv2cGoLD+3gz
fx15fx/yHDVZ1ds5AGKkUt65zaIJNOYbqlisQygz4a3kvu2NQB+/7VzRZYL2i9d5sIjR4YldKd0m
/1GU8bgH2pVXTeMQbpsgD/yLmztuZSkiLh0W5DZMeZuC/fGjwyVVMewgk42pUaPFe6adOzNfk1x7
ckm8ZwJ67iZQF709Ph2qMH4NvNZCYJAe8h8Y8BBlntMZYyPm7UIyb3HxFa6ORKhRhpfs7MVHxBkA
fZeealIVkTPSOfaAKIoqNLghNnv/UbOGG31LeSdho10N7pHNUKbajx+KuRAOOdFEp+vwxDahJhtH
dqpsIdmxF9GsNPHZBY+qmFwSzAmQPFupYXxHIZRzeX84kcbo1lopIfs5+awsGgN7W3dGPDk9jHl4
wLyFp5wUiiyON77kx+9+MUwYD0dYjUnGK7nRKzh1gy6rtBveTJ6k1dA8JcJNG0JqqmDs8gXxkiz+
uJB0fFAgtkV94wI3Imw+ID3vBmbIdCe11BD5iDF67B1kCcGjg+dGdmZKYx7PzhvcG3az+TFRmdS+
oOlUALNu0CnO39FDMXxkSc0NR/wMyKXnfq7mC8+mq3yuhroED/XEBMlne078HonL+BQExwnkRDAo
COFUVmo+aZv2vJ6y4qg4NIKzesk0lYTiTK6SMsTXdqUgZq//yvuEAoZ9fvJ9mMbe3aZWLLy8H3hV
cM49qd84OinBc0lgIbza4JHD42I3f7+E3AQmCzqIShLwXdhVRks1tZHfMvv/Ux8tOCme1XkysoYy
SgGqczrIL2+WUxQfh7nSKxHLLFll3WVUk+HAA0/qj2aSOEqi0HzUrLGadq07SDqyauWoVdEcZGGK
G5r3Ucz36R5KZjGJHpavtKLF6PkCPG4OUcQSgfwfNSvsgICahBnN+Koqd9fq8GOcSgvU+vNBi4Yo
m9kNIr89ADVTzikRIPz34iwnxhFqI1nF4ZGJATyPRYFtE5orkyxAMgyAiB2zAUS83JH1A4uZwcRd
fNGfBPxdXBloSzeuO12QBEv3qrkfJvR9Oj3G5c+oIArHqLJqx2k13GeWwdYz24nUWYHTNlRGU74O
YGWk/y2/Qi0adxNcTMNkmt3bZheOcie87DclEV47K2ZkeXVrsl85VEdmkkl/h5Ew7LXygAoAKhqS
cp9XFMsJYGj8duOZ2yfcXXlEL4ttILHrT2ke9bmGO4QQv0c/PNrfjMvQXITrlG/h4y6PkRxJhk1O
PHt3a5rKIxf0vfFbQgyLK15Y3uWipUSbuUFwgQvvx+Zy2R+FqK2KgTD0eabMRQz9AdbO1VwzKrp/
TtLhH3+9YFKkrGkRUSJDSNjmdWk79PWNZjEV/wNtsY0rewn5FUGiHyNb9h0Hhq+CHW8Jty7wYqqy
GKkb2uVhaKTOoeyJDXj25JuMIbdQ8O/Zsz5DScQJ6rlDVn9tdawzH8qk3BCL6+QqJC+mzXJoivOm
CtfglCI2i1AnayrQW+Vaa7t/5Ne++J1/wd3F7gNnTP/kqCRtklvn66ZgCpdrkhlBDIphnCKEnkgq
1eU9wHIDXW55O6ybd1ggPikT9resOhaRXmyJuFie0pVeTpGaLzLHX/wIpXpwO51dLS4xWwEeDyNO
XNp6XgWb42XPYuEiNCSpc3oo8AWU0RZQYTJrzju2q6UPKXkHhTmrZAzO+lP+AJIIBDk2ob6St+46
vg9aC3KvmcdIpLNj2TJbp28pBm1cOmrUeAjZ9UIk1V9c13wOPFFV9fdXubnJ9eA3nWRLL9sYd/O0
/M33Cw/yAawVaCePOa280/OMWbG/viMLfT78iWxOpQWo1QXlWXcZf8GoEWzDDdwRj+QzG1Wl5JyV
xZJlj+uux+c7yd0s4s7EmDgxRwJk4S3E5X5EV0rrn/EoUHZKrhbBCDtJfQw+Do5zJS2jC0dzZvEL
qjM4r1yIaqyeUDoWy6IrsIFaB+k13dunH1D9J2PeG4s+gOAWixJXBKO0Pmym8rdfUwZS7NMCd6QO
WKFQaZ18p2QeFoK806Zf/MucWbSBgwgTz9nU+4qhlRBGPc37XUgGR1yelyNfAN/922tjuOLzu/eD
9WJx2rBkL+MY4P3GqHlygByYY09RKtrYmmWic4/Tgjsy53AkgB2GhNOSXRl4HHN91JTXKMTtR8AV
cNXKt5/LGyq2TMTnoTsb6D6HPhusn/YIJrH1DK5B9litIvp8FKnyc7ABlpMdS8lFjbPlsclPE0Zy
ta6sLTSo/BbEfiC4JeLqQtRKsETyfBzpeErbTQX3DM6D2ArlVt475k2pxKtu9Jh6NAEGAyamNXZa
SqKS8yv5RBD/e30bOioK0bvJ0U6BoFb6f4f1n/oEaRydfBqTS3JtMUttsqEPdFNbzpMd0GXHC27j
xabW1iG7n9NBA1BtNDr/NBnKR5/egWgtwNSHRahcsPbN0Jt8auM9K8x99HiG1mRH8ApUdo1bwasb
12tmku3LSStq4nr3yhHXVPDKF/GxzKEnEeOcs2R3XRih41ZN8HnzzhtbtEcnoMTQzp/yCleDSU3I
+yTyvPl7L5ZxF0OOhi+ucU0asTZFGexPQa5cn7bxrQmEIipO3uezwUmJlzfTiAyI2tG7fsb4pcgw
weJTT4vUSLh3oo55GX8RBnsBNUdwTzpkJ90WSY6PxYpu6M4Klkvo6pq9xVMgT5UJGsfxC9aG4K0M
5YT86wNcg6Vydndxwg8rVLitCjVuRKSs2ROMn0dkg9InasmT2AxS3Gjnozj0FBJ8CvakheWbWuMK
v2bNm5FT+X+HZH0KMvhPq+kV+sCt7zn1sjD6Lrx5XOxVopc0aJ+Os8g75owz8JKG22ZXrgxQ4Xj/
en9ikeOQyBv0vQbNATx+xpep8+GSyLVlIyh8id5PYvqO854XoMqPZVaax2Rb7Og2Hnh5O9sOisP8
QEDRP8Sq2KeMMs1C1x2E6baqdGfk7RMisJdwDvrv7UP7hTu7nVtk8SnKC3xRNaikU/uL/ZU6SKSL
Oj8GGmD6bOcoKi1KX81voWsO1yGMiaiKlZfpxsaWaIc5jAulrV0T9VSGBy/51yHoZ4/oKZPPZkOd
ehsXdHrd5QeP1gvvq714IifuUIU4Pdux4K9bsLgtHIKzKwWvyiehOnMvNXodS+AKjGYZahSJTHYQ
ZpOf2hlfWSzhbU9JfMCg5Ijcu8jLc/3XjxRsoxNO6P64atxEsGzaKUsHxnQE7P4zXWVZolLREyhN
LJX3MTFG96n0Hz+lrKSYDDjkJ30q4FayjdSjNj4S48vORtptEVBfVryFGsJ+ITn3d5XhnULuFgfw
JoIzosYUsrdl9nyp6IjlPMLdY9VhLE7E2t8hRyThfG1WYXKBPWhLPmTIxUjOUwdb8NMML6kvX8Q1
IWNRJ/iWkOLSmTi3qBkIbRxNkrd69Qb994ZS+m1qGEe7uOf0E9ZXDq1omasXXX8qu0hU06uS2Y6D
N5pUAi/jctbFUXpx48KLWItr0DKMDJRu5N67PxnvjmCG8IGlsV6HRItFoVBUf47CLbXvWUv+MxDD
gg2zIZmqY2jcQ0nY0CTU3qfJCkEPtyJCulahUw2gJacEONNFKfVRoeqhMmqCp7PiL1chRmDGyOqw
JrSmThf/0bT9zFvxTEx34JWpIYk5kUTh/fleVZ/+EcCQbFCkyqc8a4ggera0NTksoSTAqj3DQg3t
Q4JoKNdZnDWVSyYuAghUhtxQ6P8vCpBXFCEChUM7TkrtNkmG2Njd0xjOCOs3eUW6N91CiG0ACk/R
JHsAwUPIj0lOVsqYlt0aumdRxyfOGDrhJdQQS872y4ljR0vM7V6DsKONkxcHqcMrEsGhEdhVNTA1
Gzj0xAOuJyf/4uxdOn2Sj3cZ2afuNfTTS+z/SHTz4PvNfgEcKB7x9uF0n3pC9pf9No6Roy+shMQC
vmX861ZaJSOe/5nM7rJLIUXZ61tFDG9Cp5c+DJL7vY1DyFea3yw4rK51muH+R9mEF0o8ZHfNtad0
RfZZCFd8JkpSeXKMY6YPdLsvUJWH6OV+PLMDQVneqbGeYxZzPYvsW6Eu9IgVuA7LeyIF+1XFiSBP
1qKy7IAE9BAVsKWeMnVGzsZc6WVefLwzFGW8V6/Ce3CVfJgWfk8wLmd1z/APqyGiabQFS/ToKZ3m
SQ7zLWvAqA8T+O2O9itgg1JoRwAbdpVwQaujwSI1KlQb3szxJRZJsaouaRRTjziVijqMN/dHuzr/
WhseyLlSAcD7ZQwodM8PyuCcGGhb8fK2RitSYK8YPZjIFRRWxZcwsbdQhGTtaVS9Yz9WoIJnMAJH
uQIaSpA63FnSqpxNiYMZKVwnOm0DkLz4CphwZWoo0MQ0EQQzhyEzv6+M9QuCLxcXVmufZbZgTqBA
SEp7TUJyjP5mOMCW1y1v6ZTLEsw00EA9VFybvNzU90dkjYASLPzGSfgDv74k/ZdNzgNxUV+gjFX7
uiA5ReRHe8695CUla344RRbnPEkmz8V42dntafyXmx6jTfT4dDNWA5kuiLsPfvMhVLu+/+d+AzSN
luRGhLH1252nQ/npY6PXFH4NZaWwYaGNKyeVbNCLGjlWoBSYuAFnhQmjFFmbSPvKcug5PiIo5XT9
cWfQg+BErjZWMEgHNmg/o86buGp/ewW3xHetXAjOBw1zDdkhlvzcqSXfipd7fHFSG8uiBrtU6mP/
SKR783HCVVizJmGP1tYuqmhgPRVLb85a1bfPuCbwS9VnkCgeeOZOzOssvWe1qA+DrSkNYn91JZAW
Y7uT7xvtjnv01qUJFdq50CsrwA0HOIz80+tZdSyuQqB0inpE157UGLNKwkvmNEgpZT3qmeuSdWZ6
q7gRg0xC54AzIMTXbkrmEs0RnQkcfIF+qzlmz2VhNluuv6DCshr5JrhYrZt3uVGnX+vbLbSr1LAC
6dt9vjU1puj/mnS+C4w1bbMCRRgfv+W+0F5bmo6ZHW+oOv+bbIQBEaE6hW2WQ0eU5wGBwW0N/jkg
JAOIhqlhnsoX+GNNGs4VGBSK+nBw+m5/RPGvIFaPagWMW8MJZCCSryUJibcSYRzFDTrW+Ae9ZHdq
shDFa9xa6t4gyiVg7yYdeELTstomc7LdX8ci/8Go8x69sraOvx1sJEYE4G6dhchXNML0t+0NgHwb
IahHIV+Gpk6hnBIsBGycY7WAGJFRVXmYHK1z5RtK2qfJRA1cVTIBh/nSBJvDoTkAIRWjLXcT9fVW
tfppid8Ey7deDP+QJOyFDxQLL84kp26LhBQUYGQ7EjoIRApW+VRKUC2UiXI4Bhkd8LgLi+Xy0K4W
IpixNZN2UoV0800wI+PWh6MlgTshHQJ5I3PZNi4LTBa7sCXzfvSVVkOLv3wtfUf4FALWeud8zWtF
uX+OO1iKnwtqOP4CmdG+NzOpWKfhs+HrD2UrwcxWNe+T1l+l79lG+s7ztnz2MJ9t0gNwMz1xNuHW
pyqhHPHTDOcuJm1zdGocI3Z/8sKLYwqIIM7zSVGiGtWjrvsa+Nu39VkYJq2ksYDKd/uMhTdcaj9i
rhEGi1zIsCc6D5VVAOQcJg0D3O1G0TAlP9/FQLXYmFjhoPbDkfFXgL1e6Dfw9rQKzwPTgyWYF4cx
vZuFkZ3foLzWHvCmkrP3qUNY7WcCfjVtxBOMPHP2T/xMIR8yRnKvAnK3JypPOLLo8I5yAfJYkkmt
O2THFkZ+mUEMYFnp4GMwTkuq64qRXe3myDQcN+fpvM0v6jFadxuDmfq20pKBVGwBw4WbM9qz2Q2G
eGS+ruRLpm/HO7dgF825aeIAsi+hldsqlGBvBJ1RNzdT3l/cNuMu/zfzxzMVcl0/H3KfpESf+XpX
zBGgMEIbPk7rb/JG8IZI8MSC67hGAwiPc3OVo+ggvAopkUzmZhwOG7DOZV3yZIhsa7gksM7fP/YL
ybrf2RIMdALDwDBvt+VBQnflLXi84ea4bHzUuaKcbrW6F13vFgl0QJhpfDSBps3kw62DtyPX7hX1
XpTk/ABXYiQCRgCLARdybr1v5Kkd3BqqY4d0mWn0QzLqWLYalTfAjwdtcsLix7Sk4YX4sC0Q8NZG
K+12BWdLc8CHyD7bPkEQXHu1XZDt29Y42VfbvTxRyAlFCMtCD0yGx0f6W2N9KED0KFKo+zsC/2Td
6niMtzeeW4z3SqvOI36jES4NOlaPJ55472mku+rsMYU2un3V9sm5RkqOUGRg3JeCeZoIbGOO466n
iMx+WeaPwe8BatZtLRAYi9omn1zOCxNjhlUe/8dexPHhgtYeBr3Vr69jDo9IlklN4HbYXbQ4aaqb
/SwJgyV8SRBDOk52/7udf3ZDcbHg9Dloq6iKDdcU0LIKGHx8OkGy0bVPPrwVdGThsuKKvzEwgx8w
1CsyVBMn5bUFonoNjPnAzeiGDVvRJpveAs/fsjA69NbItc6RU2CT/Vzs0THWdgvhDDJoubAWEW8Y
gei89dcYqjcWWSWy5XraaB++Ojt7Dx88WWsWxcaU6k6MObHNhnn2J7Retl21GSy3/ZwRFmCxFtyL
MhQAAZe93I6UwJjYTDRCDv/e5NMxwJpSdnuDUMlj3ZjKn483udWygYPZBBJe45s8Qrcb2Ev1qfLw
jqdn7BCFmwUwpAkCmIcPejiN2MeadVk7Hsd/AmETylWrmK5Nt6RoN0Gc/YAOB+sPcyYksbvszV+n
bEYU9u8gt1QPdWjt3SH1r36y32dFB1HJ/2Pmd2IAojMJfEog102UUqWHK15lddAG3L2WBtotOoRM
n/uKnWCKpALlVuH6E+gu4BC4QrBT0nWEm4KsCuLZI1GLJzEveGCgFT3eMlQ/OUlCTL2OffzNIQNb
4n7jTsqJWQJ8YGnKrP/IPe5MwT6ftbmHtGBGouwFBxZ9h9X5gC+W32T5PRyoRzDsXAbJv/+fFD6T
Gb+vThM+R+Doz3xDvXHbjAywd4hjK8AP8lXkPBV3s5D5LspaF2PeKGk/QXt29zfImuaaDK72wMM+
CMYXYZRRkGd+vsxuMRhP166aJjKDBqt9xyptCxbascY4Rmb8+ph0p17a8OsH8rb9SR88DUJVhGeI
8NcTi9IEzAlyJkL9E3TOyX9ePUa7X225F78pwLronokqu29SN2C8UxHr87+dkR+B+Z33TIJBVmTe
6G30wNz/gEmRA57xiFbZFlE99hetPdXUEhPbeM5YDaGvjzgdO+RmF4yeLlPUfsboUWifd/0D3Gpy
KUhLHgD4LZ/QMUbwRsiduuoltm7TJ6S8eFkZV1Q8slAuKmFt3+o8dYGx5yTc5FmR+/cQoHbN8lQV
Bcg/QrxA6UB+zX7DVZzjrRJ9+Sx49m9MyoHx6MuISv/ObTS3OvodeAUJUTuu6dZlmmTYWlDz+xr2
eRTLyPG8gX/EqlOo2immS3WK+e6g1bPdz/CzHwHqZGm+9y83AjYp498Qufc2ijbKf4h0ozxFJx+V
ANoq0ynsijtD0w5aDvPK3PyN6l0oRBvTWNjLZzOje1ptqFjin7c4WJOqxRp619oSdRwamMMQ1slB
b+HI2EeSCDH6ZD+FiS/brlF28fo5A8uRXw3i6F74OTMBKT+FLTmgXsY+5gvR90iBwp0/ub8RHYAS
xwjbuR2nkMInEpxqNBQd+nyHjtsQbHsxq73CkAWxneO84/EGYha0gv2fI4hajKrF34F6g0twYQGW
7O5usULFpiDYJmUwV2Sw0kClky1PlxC/oE9u+FqhRpPx8WE1n89vpOrpH7XByUZW08FlzQl8rM8B
Ga3rBQPTOrB7Tbea9GOq9s7KYRZYpI1WOdIPpWwQLlHOuMj83xxU8BgQMLNGVQIWOnNtFS1ih2zY
VGxl5/X/PBPbS2XVYv8d/7o97n9dmed74OhfNGFluNztgA4vHtfoI6LXkY932Tx1Ijr0+3VJe9Pg
5bbLnzPuJpRsFZlyvNJOyMCOaFoz7NyNhAD1joqQnkraj/rlzgA22wCQPv09SOD4Ecp8EhG3ea5x
09ICT/eDrH4QDnSzwl6eXXuj0tHNG8FI4reMid6/JgBM92s286NnrE9Pj8/qt7vrf9TB1E+GKjss
HJVWmsKigfauHzKRzuLvw9isSsoEeIbx4PonILve2x64saLI2HdA2p9MByNWDLVPDb2/Qb+xW7aN
OCSWLc13x5Fl7qmPHPLX19S633GlKC2snYQSeydExKWdMOjnpR/BM3BlBZPA1nPvhJbKHfIY4QgG
UyThvoaodEoyRXOGRDHqnzY0ktPwL5kMLLClrnVgLcdwjWVm5xfkfFCkwa1JxHjswQIJtBtqrjki
ROa/vQ+OZDfS1MQvQSn9Ry1H7b+uHy7F9jwDHPmA0FUesDGD9OsV2e0BbErKt53J05M9T/MNhASy
PXwsFEioPaxRydg19JbxKGXMkcDPXXkBktb/RQGn1g5nwYWDDhNzGo+IYQ7osnhMKZhTA0UFEeW+
JUe9kj4XOpDFZIxGRMY1L8jLwnelwScpIbqBYX6HX9psuomLcay8YGOZYJJtc2lE5FbenV7D19kw
OdOIHwUs6GLyznyNHdDHJUaLFekOv4V5nZoak4zcd9Rh6euDZ5a9wabKb33NVKrCI5hPAYvBEUac
0lLUqvtKw/geimj0TIwqJQez/S5a6HEwMVGU9v+LEvzCv6HjHLE/WQppiOlgYpXmFp/s4HLl0DJ0
Vyb2VKv4W6V1km9udg5xljVezRQhKiwisEq93JYuT5Gn+96yhcrxdUbsRVWGQNiK5KC7PKV99bHd
6gHH+Lq4D87N/daNeuahzH0IQqiwU9VBSxy7GO0ozcd+QzGI9ivuRuZn6s2nU10MH+xeO+EEuWRV
EmvcpLXmASm1wUntaWXvtRf9MASc0UKZRGz9jbloIwEtu+Ke2RerHKHS5mG+B9O2m8wtwzUfymAL
4y3vkn7rFBXzX5z00X7jlDKBeGeN138sV96a5IyFgsbtzpaY3Q7zoEd3DkHQUlAG/u74D8PC3w1S
jrvhShDmXrDjmRQRuU4hRkWHTrsS68jodJ86rmGCpVTr4afd60iE0fzeEvhmfJW5HWbuWctfmzYj
U6CfvbIdM/Zi/bQVsuOfmC+OB2CkXOEuoV6ai4dagtrGK1yKC3ytD1zfWSI2qhQc/tb7e2hxzrGd
WKtxWUBN2l9LYKT6nYxqNrg2ryCyHgQgAsdYEA/xDch7UvhK6v9MbgfITeWopkFxedGVIyJCP4VU
JsTXnp+D9W/MYBMmrLvGxfGkiyZMcjdUqiOhY7TlQZ951w3RBMcmMwDrteaRjrRjTvaDCO2kN4v/
/ILqx7qSxtT1G9ouSTdsgFGh8bO2Q/AcH1qobl7/8iwyXlhBkrCzKj7VFkUYp8NmHEWTCuEoghfe
BldQV99IwnaINhzqbty51dxYUFGfxVx8o6XTXOyhRw3vs7tfCkKeOyhuRigRQ6dlv90i7Eid0xNG
yeH0MhLqoow3x/QJgbBDiH0doIjVRnG2Obv3D45zNNB/6pSOps4fB/4PPk2VmGeP+sav2BVZOh09
n3zJ3h6Quf3VftcHOXeyrmZyls8dlfoO8klyaH/C8hNmIwS9RItVyTl7ncme+I4PRlbDgoZhJDCF
bsD/NzSRmxFgCGn9nlilRDi1XFGCkuZMBB+tjUwcQQc31ArzEsvPI3ZnLclMjDgt4FqCigAKGy73
d3G0pdITZlNhlEbeC+duUUk7asl2qxfEjo6If+2sfMVcojAQ9e/TL6S5OvLdsLqPUgqF0jDkJnZH
WCe7NFGO6ISzMi7WstJYgnDgp4dp61tKbVfDGh006E1ES7qjaOgmrUjmBiXZEZScvzZYIuzqjdXL
oz5FZ+pvQGwOEcwHMnmi8P6wf3zBL2vUCAyHy9sFuYCmiGgM7HbuHbaQTLCC6wRHXW5Q/jo0LlHu
ViCc/eJKYnbGCc7/pcNGsxm+iP1jso5cOHly05bHNeyyzZmdHqF3bkIu3k9Xewn563QdnSPkDlYD
1mX/FSf4yVCpiKN5IQA9CP47WQUzAnvc0HUJ4DY3KSUOLM0/pdv7WEQaRNdnB796ZXsGD5dP8od2
43r+zcbmr/VIHIl6m7uAETx6ZoiHbysZexFPx9ohlDS8P2eoDf5EcAzf75AbD94tMKu1qKKTynWz
w1EoUI/I/k5SHb8o/aL9uw72aAz1walRc98ElqFgK688bY2LtnmuvLyj0OdpJKrLBvwA0IwhV4lq
tx+/3oKQvpNChazw0EFiVDSDgpa+Z/RL/aXL6IiiQQuunQM23kNfo0Z6G57WpB3UPZg8mLPY+oY6
sBsxhAKuWonfLPWPFLtKwi/VXUmfeV2UOr//eMzr4QbOV41XkZcPpjbBCLNWDYrhVLqc9hZ1ro+H
zuvoMKn2SAaln/RKvMP1lfti64v+wP4Fpm5rq0aDxAsYsl6SOKnj4grQRYIv45sB2uvMZklVJmwF
xmw4clGf2AilEV3ZSdpTTeVwtqyyz2TrqLqed1AO65T7Hb9NdqEbGpr4K7uQSPiyQv0xgUdZD7ED
zkA6wXcPPElZ8BYb/A75vON7b/UQqRAm3xY+O4Db4pst8gRcirOq757DPIxkSP4MMPDGxj+yZyKi
x1RXyklhe/nYScRFpd4sA2g7NOp1hMj3S4fGWH3CUYvNerb1JE4UFT89kENKbVI5jguXoAwxmSDd
+V2qVN7r/8cBUiEL10zdQRmc9KVY8gmbejTb2/z6pqSn5EmdMeM2VePyHbNqBcLfT3mOepz8rh85
zXOU3dVXOi1WAeLHORdPWH0NtCL85N3uOcf68t24h5fPv95MyEIxtiNSQ7ETCwjPp/fM5L//BZsU
Olhc4CuPjgn5uzexAYWPA2imAV6Rc6nuJmcXPNMVkxXZC7QpXwZZwNzuJUaGCKvw89q0DBXu00LC
5DBgVmxegHF+K3aU5FB+mz+bbd4abIJADDU5TltvgEODgCZcillglyb791kQBdaIZXwNVK7ZAx4R
7iGalEVoOygeID6esgyBx94eQkVbRnlej0skeJ7LD7KnqBZh7lhaR1WUMxuVLNkFIgOjNsfwkxqs
url6vGjEberO7RFMeCBuSeQhxd3Q1u3pIXtCMRhCKJ3FaM/umzokcnTRNbEMxEovzfnU2afEpecO
4rvkoNGbNUVoTREXWpewHE0tvMFaeFrMs0aZRJdmkCTmizllODa33e/J5izkjC36mIYMh/RoI/Qo
1qpqaPErHAjUuibi3p+skmEP9vKOzTfyZA/xUvzarnh7eKhsPCuZyHrJqaCaA8ke0EnEOH6O2+bf
PczI9592gJeMEwsrn6DDqs2fmCFBDZPnHfLpquzufpUYaunG3+vrW1cDxoWwG0m/GSM7xDFKcNpt
EdnvLH2RuFMBKo/V0oFlh/gK6x2pDcEEwUYEtoUIhGGNrtYgAzxddOBVeJ3oocXcx4BlSllvjgxs
0YRkuwXdPG5nPW/jQhwIoyqhtKK5/i679OPz/JJtO/Kvlc0xosEgUdPKCgxrd2hj7rnCephW9CnC
RDTcnE7iLDH85NjmqXTXG0Mbrrc5iQqQpfksqAYCqRoH2s/Y1FmTbCXRCQ+vggt0zn08ART3xSvy
xIv2NOXI9HsXrz4NMrqFTfhL+9QFrhi5Jmw9bKtdL+RmGLs8U1Ha5gkyRDb+cnecTHp4nA6n+esW
U8PwE53uNgas6jclQhqnrVwDivXFip+pptYIljoW/QiW3gHEwK7KITf70GRGeEz6u4Kz0oLHtZRc
T1Qcm3SqYtJzctlJxNuirMZqKFey/yhwfezAEduJWqHSiIPEpU/uoboJpbPciIeZVHfMGiIXoVHb
J35LuEb6QdjkLszd0td7Lrfe8hC2A82/zPUtQgm29iszf6q04WEBclR7lqmLhqG4jzXM766+Gq+i
sbjh5Y44RLqv2psdQ9lKkBiU8Fy84MOLX7R57/MZzx8xme0S2i0hKizoyiB+4TcB/iPugnsKImxI
1Y7DHcDTWO975sTSUBDVp0id7a3muELpkgH4hM3dPX1Xg5DQsADJtvZt7x7p94fI3NMlySE1NXen
Tp2KuUHGPEdl1uPo6ofmn2wugcaSKEmQbrGuYufq6ZlMYHueEHeliJCM9UF0avwVwKzGjUdBF2/q
Y36xVw+EE9Cl2SiejXLzF82G4VeY+qvolPiwbDeQz7aYyZrt/ZfCelz/1q4lwkwhAreg7S/yQia+
ukJjQYoku8zC5v+EQVDYmOHIkgOe1TDRQG3UG8pDkfTKHXwel4nC25iljMyoE9EswwNVWW4b1pla
64LZwfs3H8HCtbii9ZK2Iuiebdohy+TPDqKQ9BXtQPb7LSU78zJ+xnYMLB5whYY1g5pQGdyATsjc
/cgLvSSS0frlYF6znHGRqxHWSDscTUHm0hcfHubKDHZ04jUFJ+rZKQLkRHgPd2evwV4Ba1TT1xN7
6GIFoiQL+8bB3piML9+MczvZQiSGb1+RCWhYi7pM5Jlo/7Z4HtzrZ1WApbCU/hB0OgGy0FINfqSZ
y13tkgejxiO3JywTYOj9ZRk6b7BlznVtfOXBJymk28h3Gpvp5PeykLr+cuuMPeNZsi8dZwwvFIbs
NHAQZRlpcju+5TkDWCjxUarShF4A1y28T2QeyzXjg+hYLXqAkgdqFC6prG4ltTFgCMGbKNNkIX7d
7F5YwennTQIk9bW6h7oMpAU5U3BdJgrR1Gy4iuc/2O5+dQ2yi/+AwZSnlGwxO8XkolfwM6e/ACxt
0lXNH+pw1nHO3o2woKSEcct9vGKtEBmtMgLByB42MElrlOrmLv2eOiV8OofSUslh/HXHBNk4DgMy
2QmYVpxqLeJcLI7zBtFK2TmJ/++SBon5SdFLCkbeBnDhlW3RtAQJnjDkLk2WchmteE9I5yaRhH9t
FcyB3JcqxcdagJk9/VGKosqv+05oPd8ZBapuS/yTNq4sH4k2I2tQ0ybU7s+X15qJJAJt7treO16R
v8vQHlKu0vYiVmjj08bOXTMdWL5xcnTPMeUTE0hRwXWgGh1m9jMqQJJaqnvF6Z9bypqebZQ+XRX4
QZcL6rd3SCIyIAFhBBZMMWmZAVTy2JfoxNrP1Q8Re3u6paTgR59xzGku84u31tYPLY3zMmILSfWN
GyjNQvFiPfum4iTAoBL56k/lp+055S6GMrv/vGL5CofGnVZW4nUROcoeyaayQ3yAXbdmg9sum2GR
XC6eY5h1exvztsfKjDeIxRBs7KQdsH/MsWInZt84Y0PxTz9wknq/24522q0RhGV94zJLfST6HIRH
JYYNPm+bIN80AezPbUhPPlqQ0fif1EoApEn2gPkTRuKzIeQ7rHE46Bz80uW+1i2F9Te/2+HWRlah
wJf1/5fdSMINfLXFeRwljB7wlmXAoq7sEsAeO+/2fGtTLRxNxTC2qfa5Ui+KsRdOrhcJGeQ2sBMf
6d6Pl93nFMNVmCJHBBDInsNT97Uhpy8fVp8cmanV1KATgVNDmISkPgo7F1KfSnTvHtTAA6hUSMjF
Nqk+aBv5B0yyxrfJCkVqjnfR5mfjR6gS/aS4jFNWPTWHsEurQ/CAYjJA8gWgyzX6nwOD4EyqMfd2
y6zx0fEaiOK8r2/JVc/pP+y2uYp5hlch9Pegr7Q1i+R78eczBW9XQ2jbz5l9LgDOhN7OUuL296o+
KojIaConeIFwITGM0CYCsus8GcQsdjGL+hLj90Wfs66/cKyLwqCnImP3qPhDVndq6YtaZBfuSt2I
mDXKOXETAC0+p0byzdfILxa1IYHwOQz5HagOKskvlpyET831hPZ3fFRR4Ut2rAA5RJ9qOIMbHlcK
yIirUJCvM5E7D8EBRTmXVTUrFmd27G15uH1r7wUvmAD6OeNAO/oNajLsg8jf+pUdVpHSgfEnMSbt
9fA8jw6X/KYS55b6rp/rIUVDQKCpezzNtA8ux/OymRDiVy1/P8jVxUicS6pVxeMCBGxxFnf9og5l
SJ/wBVPB3KW0c+CefZiAbgMB2Vtq1ILybnOx1lziE0AnEgrmmpLNVVr5lCgPNLqbB3O48U/TylSe
ClSIwTE/3FGvVHrkchNjP/AutqqnxpY1Ze4nVjEt9lDFo4ZO93RQRmEG/45KqpGUfJDErMomwAdH
IbPjdpmpE0CAOTRn7m/+5hUgQDqTC1HeXzjDrIt1gBTQIGgN2A5wSVyXegyqhsubUZ3nCxRXF9rY
iyGhOraUFPY3sYkFGmOpuz8gfgH0aaGKHBZN+2DCWTq7jo4XRUPlYj94SeM5k4Ys1StGn9ZHRccc
UR/7mHS9RrkNzzNVd/1ErrFfdX2yxQ/Aa3Ehz5sKM9NU3G3oDWXpyZxt/iA1KUx8tbbMJITsZpQ5
e4Ty+1cDnr2zELwZOaG97JNckyEIAe9kAeHcgTxO6tdKXHp8q1QWiSaK8etosADysZRV2jUNj4kY
mOnc7Kubucm4HhtmlCQS7boj456DSsw364t9m9jkEdLo3MqVlRVElILHYtTweahtk6OLmSDLNdnF
OcepPZl8kjR7owlq2cQjXzz6jhx9lJz6EqePVzK38r7Nzcog8fibtupumPHFsbsly5GqQ2e0Jm9v
hG3qkA8gFNQoERITeN2supgAclGwg13FRAPy380xjBU4BMiRbHzAI7a4WcLoQROozvGwiQL0uihJ
ukBzKtxUJNu0DXwX9TGTU75xoICJzLOagffFOlD7lJrrWNFjq8xjoTUnxBkYKtipJk87AMWCypPg
eMQZfpZijoTUfuObWfySpVvI8GfK3/fQ3zPU1z1W0phBQAu2VVo77UZa9slMmYsXyK2424fCCs9p
lFcnB+5ex6ahzmS6rcOYG8BdG4d+zB3DoQHMzYCXTZ2/DH+5icXjPaaRvy+1VN0+wSW4NmfveKip
n/OlekQNg9kVaK0wcL6umMPViTTgzMiIvjK2LI+87XtWITgHiz9y/JS8iXcq8+J525vNVLBKop6J
+axEvvXg3VwqSo2CtYA9zUFyf1ELeevS8qAxGkhsIAQWX7xGQ+vR1yeds+Fb5AS5Rjm/Jlxc7P9b
/f7ih+3MWgwOcgfBB0d+BvsKt/NZ0sE221oiFScOYX7KNW6knp2AIxJ2MZKU5sGgKgtTTvq102Ic
TzVc71UNFA6uKBafAt4bHS/2qa1SLee5OiUO3Ba+pwIyIlMCP+1c2505WLwVWyciQgl6mqOtw9BT
ky65gLX5H5sfpRqIeXS6yv37uo4iGf86UA0gNpYnewL9IjM2JQHJ0swUqtHQBx1GDgUT9XAcL43o
2IXOvk7GRr+XZGIotPqkFKkOk8vI1wiCJN3tYcRycBEa1h4h+WKOUJoqMgdiKOF2itg588QCviN5
cAdadkPADEpAFNOJA7Kvx2527/N6dJTGkfdLxcUUxZP8g0Wo55rk+0MPdAKuVUwTs0jgrd3d+Fw1
oIne5d7o3iSHueACWcdQdl6DYPkLbyiaAjqkMLK9oqr94RmL6hPV8WiBz3QwuRhBDauMP5i+sWU9
j9Vc9fbYfnH4uh4247RnKZxv1s9UOiNX07h6vBBLQVJ3Vk8V+O9/RD7K8WD8qjBdHQtrsxGV/rbO
602ErCIRXGYAhdL5SiePTz+249YmuUnr/O5JM4l1U8le6D3Gj6n7z4dMEf3yYuwcthqUrBZhBGxE
98VP52InBeYWubjFKty+CgJNItoKufQWnqlAaZp8oOFvFbthUQjDpZeSsX60CyN23aF+hfqOFged
UDpPJQrlzWvHzQ2a/qYuWjpd3M/W+a4xc1u1jX+52d4/e80AeOoj0BarUHdgjGdutBSUGPqB6sXv
Mg68iVcDAmmzavodrvKRWcBb+WomlcnLT+jeX7M5YhX7/6zgYWmuMJstWO/+uZ8P9WXBkh405vu8
FyU0dfyDXZU+m6j5zM7NPbKJZFGJM/9ypyAH9JWi26jx2m1JVobaeI6L++HkjRCvTotwZBya2dJj
Jw4Aa9b7JoJFnIdBIppX3XYh+JZOeJkpxR2G1X7+tOBVHzJHcxyNAaqajYCSVDSKmF3G5L498UKs
HtyG3MaLOZOpWJ0OKV2b+JMabGI3rTrZFfoHPGqQSbWrHAHDJDsmiE825MAFGCJhVTgetj8aWtbA
L6F1+1jLvXQoqAbeH6UnUX/we9yyPQcPrvQjAXWTnHplSVmABUNWvFNao8mQLy+4GylwF9X5kebR
3gRx75Lx74LBYETxRov4trlpjhI4VFcgOqVXlPRGtACOh8q3jvkO9l41cQVrONRAn1o13diPIa4W
R5N/SZaJ7JvNx5bXYv4ll6sSoXKCc9PIusbJVKyzJwooQULVQCY9tgoNduw9axGKA4Cy+jOkJGiO
0woI5Sai64vTxK3cljSbsuKFIlM50RwXwultYxsKKxzU+m7DcRbtc0/yaDJzjOpjpTgeWxJgSGFp
C9XV/B+doKlHwF8kl+B4wwh9rrGwMmi5XaKZQNrpN+2nS/uK6GATwRYyNLRLL1gK9uyS9SadTL0s
bKnKXNsWsD8fsTwTQyt/HmUSKuQ2F/thEGhwrhWsDb35WBP/nso8lalOKCgGXTZUnpMrgoaDgrcg
+qfVeV0W3xxZQhGJSTnECp17rARpiEDjp17SvMOR+F5VGWPSqE42upkQddxzQ8ls0EgHZE7scPh8
khNe811A6YwtsQFAUjfJt/XR/yDKpnUyjilXDffS5FdTqem6X+vjyiNRh0xQFexcKR6ooIwJkoK/
/N4PaAjGcxupCPXt8NWF52a5gJVNBF7jhcQpbSXHxYC84tacFtfdQuEF7tfqRe3vpzlZrd+BU3NE
+gFjrtWRK2Zq3124dr+WemBMu89+wy/TQqHmkHgi/TBZToSceu7f2dQBEQXO0LUMBFtKpF7IHYVb
3306/+UQh0i7ApYaZ/zIOg1WE1nzQG0T/1rJ8sOaVvR7UdGxzXMf+peytdvEpJshW8HMdc9Zk3Gr
oIl+gQ4mVm8xLs6yemGbK1tlbOiQh18Pa2pO3CU01w2d/vd/5W6izoBjfZO5yfUnUEsW28q7w7mg
hrZ76sGOomsVCedGObaO1sAM133n30CZW0EMDP0fg1u5lH0YjItGDXxzNa53w7JuCpB9VAwHs/IG
GEh3+vrTTWW90WjrPdUWSsYm1Hjr2ph09cejIqzibi2TUo4EvTyiaeiglE8bntoChOquIHkW7/W/
CWHDijZT1tWf1+ylWrjA6FIrv8TW9FGtjtQaOUXTn+wYUrqpW1SIZGhXLxFk79/SEorY4mt4fHdn
o3ULEaaJqDim0O8D66Se/sCkgMSr8eydIViiyUvskoNoA0TO1TanNPrVUhNvXVInKBJ0/t4AP1Uo
Rxq1iGwjWrVvkzSMPOvaJhSimEGvDeLo3U8AZunoAT87SCl4bv9whL88p/BQPVTnLUvInx0uSrHD
SMu9AkIJ+dIw5S38RpEEV/0wDpQL6haj0jy4iuHIm+GMzarLozvh6q8k7qbs8iw9jRqickgRYTQU
pRrU1rBkTRX/ToGeolHmJxQLsXA3pBL45KsL9vqQzF+/Ng2TqjJbOe3sqpqN/v4ygMSgG+N69MVW
WkQ5rLYH0GYMX6cX2jIuA+UPWXrncBsDzurgj+eVsJnJkVOawu9uH/Le5yCyzBKOy4Vrz6ePbeON
Eos7TVOpZkNFW97iE6cO6slYGFfONFIs8MwXFvAI/7GB1vVc4UnhSrvsczaXaWw3AZ/Y4k9jTMD7
CAWlkIxxJWAd5S7FfIyNE4aszpMYg7sS59O2encW5g62aHzob6LZHbD+POugRyhf5iACevnhEAhW
Xti4hF+eJzN+zrugk2XKR2Daakq4p8tJCFLs4xULvv5fbOZg2CSVHUH3y1IjBRdKCMSflX2/KE4z
VbBdimwoRsEXY0Y0uqWaqgFLA5OtS4K5mc6pZMfrGNXM2Gc++RNMxFAtK7LhBKblX6GPytL5ZjBp
SeFpzsHHHpmOyCQuPi9FRTz8vQ36Z7wRSO3vrECj5XjbvOh1+0M61Ovw5e3DPu2jdWbZani4vVhX
tsJTQjvdA2Qje0/miz5fNSOyt61cP5RtjGZ2e6wRK499213xHSz/m5Y7nsaCm0sceerzLXQrXtcN
0M6ZMCaQ5jAgoixFOTmjL2NoAdyECuowVMIiLOB/jgbP3acSOp9Fz8w9wsdzm/mewlfIZRv2yDSx
+bWuZM5+d1jAbXHU5Xy9LrkE/ZwG0dhq97ZOu65RcRoD5Xahsar3UsyVc/AuOZUDzbluDfQnFTZy
49V2kbc/k53g8/Dav8BJ3v0T01/4F/d82PMF/GWwjQZVe59BoV9NqCp3AQhKhkXBEszJBcc8pkJC
+kaQWjcg4f9Fa7T544XvdKNEHM0RxnfOGwb0LViyqRRTIJyUI9xgyw8aG8Eadl9buOhp2r69S5CD
vf+rA0gIaP3aFLPiNviQaIxFkemez/vQv/JLBcnC9Wq68IcC3dF99x6kmroiE+03kMQgG8ncp9Ch
9eo9zvUKAFwO2MSP3BoPLb1xS5NDt6ebpowdKFh8Llt6gZr+sDWZeQRx6z3jU+fWSSHIfb3Zy4nV
EJp19RsjqbuC2+mdrf0cOY8nNl8IQc4kh0s0BHtBT7dm22fe9si2WL3r4SykkgYAdKOAUJUrYW0j
nLbQaVqrkSIIuVkoqFlxFbhvGszzNa4bEp4y7jzODm2/Qs1TOSop0IDTioLO8vkKCL8PGr5H9kDz
k4H5601DSrNj2VQZiR+EZOVCkqqo2ilj4C0cnpLKVvUyMmC9Nd/a+Q6R//NuQ4Pg/j7kcgmqbDWr
G7vhZZ9hv+qymAKncA/3ney80fVa0iWVMf0AMVT46NZoyvtQV1Ukm0IzeuGe2zuv1C42u0Un7fBT
ZlU1sEyTivHjx2MWWZ6awtuWCU2rfpS/6DeMekktq8TSkK2G6P0wxyaNUgSE47MwwL7wHKZqoM6X
H4gHkczaBFlsyBPo2xJZWwxKo5vwPrDsKgrcEfHYviv/llQqvE4UYAxcGC5WzNxGxYhg1JkPdE1U
krseCv39Q0thIbz6OFaGtY5DIfBgq0u4eC80hXnWU4sCrpc68oTkNeEYOeyNSzzp+BNv6c6g9u4d
50lhHr09c2cj/WKlTLJ6GGk5314nv2Ah4oRfOnpKy8Fd+Yp541G1LOQKO7+VnYUXfrZ+jzFs/aq2
BawuGpewzVzl7wnyXlC9RwIhPT0iFZH0gSkZ5uQZEhizJiSU0DXH4KjcxZoaU6lvYQMX8XT/XXM3
jfK1s9xA5EYd4h2Upp2ywNyyz3nAVJeHg2sNOIVFkKQUATCO/v0fNnI75msRL+lReCaUYHvyU+mJ
y7HjPzMZ1wfCw4mG83hwm5RODKAGXhl6cW97usJSiiY3LeB17W9Kl/6SeAqYrC26MhiZavsqzI9/
kIkjFQnv6fBfGAhhDpHSLpau2eKzGVL0bLA8aEF2UoGBQLhVS7x7NvcNcIB8OQdL25Sh8ravUeKP
WbfIfU6gwJ/lb8N/0ZmtHXt4yXmG54QRzoriSBUli767vXkwulci/XUvSDuKfx7ti3XiVIYkrNT5
VBH4dlF+0SFZQwE26dSQrFC4VeXOH8rf95NZLF9rv3XzmgCVH3GqJRjTOeIeoovXIfOmjZbdEj6x
P53Kq1u4udusId+uErAZGltRnIF4dOzBNMh+uvUyDfcsiChd3eMoM/L+KPylgYFACm5gZNOf+9sa
Bdgjg+fOa8Kmu6eNTJ9gdoVcJxMcfZ0Q3bTzrI0N2kxcvlQCvT5Ls4Nwik2KmrhgDjFzdKt/YOJ6
AygKnCJV/sSRQgPZ79tmvymOblkwUqyAvPk18cq7q4Bea8l1YHeGRv5dpZ929jdAQUaNvOokcwDa
jpGUDJAA/I6UBxSFjoYt/yFNWLrxRjdrVyRIaltIwdV6CR0ycSmuu3kWIWNVpGHu3Ot1Z7f0O5+B
WCl7+PiOmW8FPheu8N5ko5jXLtx6sBuzHk5Oj7KbK1KsdTke2a1DLetOAFHYVPgnsdhEsRiUzuqZ
4x60GrQ84eNfLO6HSrbOnsYX0MxQLgCu326QMBqtXR5TVkkURpQIQidUoSeYqR0LcdRaLEZUF09n
LSeB798ZLWm9ArVVnkXL3JwT538HAn7DgciU46B2eDpWsPR2j4qVQwLzAGC8oduCaEoPPGzzJZqP
kb5OywrT7RIqrXO6Tps9dinRB3MvlOh/pKE4rqSaVtfiaZHgvhcBgyp/pSLgZsgLesqf1Yu0ocgB
/38evNucu0ajEeY1NCEEA26mnKsr7qr7FnCMK4/wRNneRVLl1FcoiCdFVD5UnDHiDXSM5/P5RUTq
CCuV0ARXaCLfrn/eguZiB5ie/S/2Q/fiwivBHFxOqz70qH1iSushlRoz4uTGbdRkNr6O0eGEHd10
HuqllYkxxS3+gCaFaJrZS9L1hG2MNUYha9MSeGkgGZ8iPe66qt+0JG+1lKh6k1bf8qjXCR4DLdpk
Wy39IrKOSTHdYb+OcxElDCaNC8xWl5njps9MTNPEqO+8KmOHV9ngcQ3n4916n+RW4uD3DvK0QncF
ElmhkdJLzjuB0CNIQeY6P74cCw27DKFw1PgHri7RJW6QD74dS6ZnVFFQbGJdsn8IsMc1uUCbNPPf
wHgGyW7dlPAEsgD3BXyoxx6qo3piU3PfXExYsra54IsIszkr/p08R5KIhE0kt5ebApX13OYNHdxQ
d8jv6Z77DrNjhe9cx6bMGWtqoMCjwZ3pSa78QZHF1afvgZpFFWr3Yxuj1ZqN2KLGn3axb0tBz/Xq
YLp9p7wW9l91fqJpNqUyuTI1o7vLdZaRnXmEf870/vokmDdym9rOmgyJnWEtXyuyX5Yc6Dw4zFyB
gCN/FkgwFomfpivYxBP1Hb3phuqtD6G+ur2pe10pffl3KE+YB5XVJSd8MB09uw7F0YVrNUM8RZfm
LW2pTHkUyXMc/wEdYnqG5HXx4zbbur4FVYRLQCZv4kZcRQKkjBvyChe2p3ehl7mprHJnm9QbUUx3
QAmE92RpbB0XdcT8+L5X+M5Pl4p+kK9N3Dzb5t4/HLg++GiSyAUWS+hsP0b5zw4XWrG4zRuBFJ+k
YZnPCzkdwU49YcjUSbRi+/SGpTgZ69XkC0A9jrkMoXmfAP4l39o1mA6FpyZvF5iJIJh4XWdYyLAq
U8/txymg+o4eD7v/wusdZGqBC2/YnvlTGhN6pKkmsov9lMrgqu1CwiBM4Tc9TVxNoQzoUVkvoO8U
iUDn/JGb8UTSFtbL8Rvc7VAI2cssLnbRRWN7JZWh4YqkOdMPPxIJaAvEvlacELFuhBHX/GUboD31
2KMzm784Jkhabr8imqfZ2wilmTg3ezVi9magrRvOa8jU0yEV881Stfu7HiNbRzjo98hjZ9tJDiIa
2wiH66G3FxpYcYosX8g24p6ZUOAQdYr3zxCtsmTJP2Uv9IOZRRRWKDopW/ottq3+JUJqI0PxIM1Y
3S8p80sBLo1amdwv8ja0LONFKKqMjLNa/peym0wKmH5ryftqXxdJuC3xC0YWLHt/8sF24kbkmoIj
xp1hYJESAuXUNNW9odsYSnxRcn/uKFxFgWrNuLPvrIap7FvyOzuiVSJvP+x6GAjCc5oYITqSOE4a
ba7pHSeiC3VAGVLQ0LuECQuVHmxhnSx/Re2G0ifFuoRXPH2s1o6yAh+bxJJLrD9kNhaJL53C+iYX
CQRuk3Ed8+7fx+gIvzm/+4gXc73PRZeukyCCDXN9MHxVjm16A983PHl2IPw+d6IHUMeda09D+vrV
Zitbe6Jq4quetwdXb46/yH71r4N05Ne+4L9tk4uDReUIVlQWfeJt5dA0fQCLPsHpOlxiNUb5dukp
ahUYkhvvYx0xH3+tT4PP24CVghnS5OQMjczQKJVqrMhVK2NYpkVhBbHpiCG4rxlXEsyLXCZCSuOx
PNhCqp7R0w1sR/L6yjtFzJw4W/ogauEn/jMjgOjVvoC4+4Op76PQlPjeDUwxFXwmAZT0+JdO4Qm5
6TMjC6OlrGL/vTdZAnBRk8hV5AuFNuM4PoM7tL9Q8eLzieS9vP7KAQnznHgGk0/Z/+upqCOxzveO
Vt+pQm2x/q+IFpqzvlZgUSxhNZW+EGjRl+IGyhNyZDfbS7xTeUnCHE6UVoTwtKTZXfUNRT5pIMeE
gzQVJac51zd0BfDCl6kEAbFG2854eLRtVo5lWBCMWLDxaTz/vpss3Rx35JO3cTCeh3zxDFbdzl57
r1ewt2Ymj9t9vpPxqr6gs9w+0kZCW+T+1TiQYSUtIz6UiM4+SK973UXLV0TQ3HVRfRZ6I+x/RVys
Tb8c2Q8X45qOaRy1oVE4E5AUYGc9OID/BPLUQroGZvQ1A6TI8NR/Wxs9EZeI4sIxV3Xoudfz+MpC
GgtlxYY6dCSaJpE+S/IrctYAJQRRRlwNywBeGPCKZT2CnXoR08uSqNcIiamFNycH/djOqjdvKhqA
3pMMvPOAiSCBpzqu24quhGKp6jLJZshqHgQZlJ1y2IneI2cIpwQMN96A6kAS9OkxEuwNSg3GhcSm
6rZXVjG00gf1AZA1uOb89KHei6lGGQ8R3LIfJVCjx2jP0RipmnpHBIA7qX7Wsw3ui19DGLVy2lGa
sV6+pkREzf/zZQ5KZL6EJ+7LYaCYM6cCtm8DbFht7UD98TqMfWTQFQoNWFFKOytf1HHFedzJpFDb
ILrxq5We43fOBvJ1xptt8ckj1Vq/74S9JwdQErEenchi1unKnCAKlr4jFpzBp1cYTIQ3PrKv6GZK
iL+j0+zJQRj9Wik/vUJfCnyiKmsRDFJUzh8Y+D25K65NF7S8qSw1KUPngV4Rfkg45o7oO761d/NB
zowF91OYFmyNmspmqsjIEK13RoMEr5IVQeJLpFLGIhdTG7MEricV/BHUVHXERUURmj+K/m4/UTMm
vhlyucfmQ6zbiPV5ZaDIJng0I3gwoaFteYe6G33zRvqtr21VMWcFkCLlMlzTXaLPcXXK65PcdP+g
Yi56rCO4vrRxieWZvsWJzo912uO0YxzRKEl4KbLaPu3QISTUnC3ukzTXH9qm6UeXMAHWKEl9TKme
2Lv7iRoZ1B1RAjySGFyKD/OQySQxpO5hw+yA3GEyV2I/Li1x1COLK1hSol9YnvjFFxxCBDHaHW4m
k/MQE8NkT08sphFybtrhraanGGTl9sEhzK536xpnj2mR36htwEes3cT2dIvWUuTsG7cETHHfZmL1
JejOUQ2IEAmDbhsX5/sJ7jPIFSU2ogqdr3W861baVQT9QCc0YLq0J0a6GXhJ700ovf+vnD0nS73g
RPLWBCC+irutzswnot8LuZPotm21JLSHoYEto8iJbvjDcvi4hqq0Z5fhTCTfwABYCCDmXku1Lapo
/rmolLpBRhnlv5ZcJ0MrCEVy2qcyFRmIWl0inQmLMIcCdrcgVpon9fBAtVnXJEVoVCGb4HUehjJl
oqEM/AQHHW8vs90HziSc5iab/S6jMAw/Eo8m4+h9d5PaqN7s91c53iAgEyEiHQfBMXkR4m1gV+C1
Pz+g7Bd2ASpNHI5aAAl2b61H6EX6BngpDGQ29To2MdQbnpaKpsaZj2fPWkhBn9R5dDHz3Nj9qxTP
Vsvg6irTVaTtopukxm5khXSesdl8u1wxYofwvSMJEd+sEqMETWUvnJuFO80Ig1PwfZ8bcjThcz1m
s8ljK8Zm6glAUJfVY2SiTpepBWk1Hpm20JmokcSSA9vulehh6hyP0TWPnYTfvrPPtjLtuN1m8o59
gtHcQbwX6+YTUpDLK335srm9jz1hm2+TPi590VadH+ErqdHeh/Qns2x0G6mQMUtLm+Zr6OUKPtJs
mfQRDZ7wVRyxgsXZ/7wv4bxwhOTKnnFjCaknrRrw0rVZok9NkfxTUTIFQdghnp4k4g2C8d0yfF7F
Yyh5ZPVIYYZ3nQ+vmwaOG2lAKJLR4SOKAZIOdTqIW5nVPc8socBQLcsnqQkhqITjc4C7ZWyrk26o
AnmkVhoW6nJHGK4zEBXwKQYLbAnjxaMDR7M3yqNoXVIg10eEZocZM8uiN1B6sIVUMbI0gFgwsIOP
sluJXyZIZ1tXFb/wIs9xxST8+F2Hhb8KMdSHcdStRkASsVpWLH94ZwRLaKfpedtPKFxbNVZiTf1u
Zulkb9NnlPo8geuOQmKnTT7PhAR1R8jWqMzBD/zMbnfueqmZWVf+fa5frolF/lF3P0PyCZMSovkn
0lY/TFcFfM2EWlFhZoKWpzd91DjD5wX2iTln1DINl36juEnM188NlihZUESp40MGZgtey6dysr3f
vbnURzWdl/EjrRkmTc1bNVgq9Tjob18HlhScF3YlhcmF0/CL2VlTsWhNKNwGMUKTs30kcSEc8vQC
+g1PER89tjlE5SwO00bV+Cq7B39xz+OgwyVPpTbVZUxLbBeHW/AEJUPR4A9njkcAevoAe6m23Xpz
g+ybK5CMBON4jZiUvK27xH1EDWqCB+/RVA6KIKD4eHThyIhLFGRKYEPHgELiJwXBfMwskVsrn1Az
VsMzeAEwRTH2rh/MvqofCMyAAw0XjD8whkD6NnCZ3TFeA86uOzbf1QfQZq8uohQqhr8a3AE2FUIn
8br0ukS5g8BernW6sWBGqvzBb/M1nj/FGKU1yDPJaQIpk7oxVo0OOt6+JfoOw+ekZLvvEdNg7n5z
Z13UOlda55fHQAoAxE456en4DMXUB3jP1zbC2gOfz8HKVvQPNwPidhCQ/Pwalh78be7pvk6XliMS
gHPoBUIckXKsv/uiUOWEvHn3WfBziNEBmkPTleTqTHWCpzAgDtiNT+Y7oShP/q2RtBvJX5k1fJ9v
OauwOBxIWCFeykTt02cG57nGhL0/WLw0ja7lrFuYe4VZMUjaV6b4UyNJDnOlbNMc8o6elOzT8YYi
xdmbmRrn0xJpNd562oZUImq6HKDQ6c8bF62l8nCfuJv2YDaspUVztvwi6/lGqYD4mytO6Qkuziam
ip38bLu3mdsm3QcA+buTyKPR66CSzHdwgklchVbWBmGi4SqPwmOSCjlXnqUuXVys48jQvZMxdBEm
4+3gs1Ca4JjtqVO50Lvza3ucZOiHP1m/wfyAS9UZPX79sj1mHxv2qZiJsVHGwlcyXcosp/y9L7f9
BPmegdu3MIRzv3p2qwW1Ydwf/YvcqtEauaCVdGv1gAQACDKVALcneP7l7HD/VRLBwafXHX7+XQWJ
hHh/00ZXenwMptGjb9EwWRjTDqEftBjCxF6JDrjEaxjmOEuP18H9SiUyYmKE0v3GphkErF0gN3kW
52VbqcBO1U831xUs11EXxmtydaZ715EDVr0GJp+l2igg3ednxDJosMVpBSJwlpCDnPqjUskjZmg1
bpRpvZroK7PxmHrF6hZwoAGkZJXjuUnz0GrWXi2t09oKPM89dbb6ujIu1iXYM5GDaV1Q6wuCMErt
Oa4HYiWd6W7uDCtsv119lMEtnSxA+VaT4w4takAXfsAJqz6IrBM/XA6zkTwJ6PmxZ522s1U6iBU9
oXYGuwAvE5omDSlDnLMY8s9on0Q1vGXGXIbnhEOm0YfgU1KasMetBwEk163/nGR3tzVm0hMgSOm3
HbVbmzE79WhwhYMRM6qIl6pox45II1af8QZb5mahDzZ5OagXb99y8o9aBZS+4VUfdVHb6n8Q+qmz
TNMGSDKALtl9SzvoG6Hx9/1kLJ0BFu8/tdG4weI4UCNpzq476E3ppFFZqu/1Gk/EYT6/9QOcT/mF
GsbWbKHnza7DwWPKTBSxySGZZtXHrlmrF82q0r1wROZyB5cicwjez9Pv7DK48KeO88My4ilZ1VlQ
7bCYjqSulC3jJ1x4ML++2QPv+mv63I0z4Api3wQ9vUXbI2ecmNT6MhoMC39qGGkhstzR08o2SuCA
LrxUkGlyV2l+8DkW/el9j1Hi467E5tQEv0m69gOKOQAkfSytSofjAw2rS5StMYoSjxfwlQKcYGzz
hfrlsB9QO+StPrR4V8DaASHEw5f5l0ujY6+trhukIOu3pqZRFS4ezDj02+jXTmKTUTTn2LLRgVTj
5YHY+0tOJeAULK9Zi7pqoZeV8M4U8tXAnfGlvCDOcp0YWxZrnosaMADYSP2Q49tjh8JUYo25dgID
fX3quJUc8qnEvL1l5e7MttQLmWXiNik0l3jyF9ne0q2pNnYQeTuryhyYQCIuVAPEk2J6BuQHKPd2
VGES6M+eME52+qL0u72pNn+WPCsXJZA3wBuyw8anZeNXsQDbXNVoH3M2CeY8AVEA9WbZLghaPaEh
ctwtCs/f4GiOHZIpERv4Mae0l5OEsTGlCJMQ6t3RZYEeTWaTQ6lFaEX5J28uuNFD+wO71knxdkm8
3oNT1u8nr73aIpvz/rwOnTblt7b4lKoGs59r09EsT9pLz/5XgspYwa9KI9GdpofA62Xt2jLn4cVn
s7Gdq8m9a1PXr+cDBFgtktV3Mc2Xr9sEOVBFj85CBsMkpuLEcrHG5FTqHbKL008aTj0laM+Exu7g
nIW7qy/sHe7cPriiSgEuBTg40MgG68W8MWth5W/749jIPjIyPU9hGG1rcYgh0vszJPIJCq8763Mn
oP5Cja0PMA0wsou8GLi8f96YDzrKXSNJTmWrzU2Xc1PmUHDfn7pq327JtSd55NEvEGHUzolgb4Kz
iCCD00n3jInPMdW1Zprwh2yecP6XDz278OwC8bPUvj5P82w2448hbA2wjYA6O+ofjySUSxdoNXl5
zv+0BZ8B5T1bdgmE9PhH4x5tUJpwEkeaaxeUqfaRzlqVQ7Ad88q5ajQrNmccJIxSoQ7raq9bgg0x
xsJK1chS82fOfmqc57PuioNBp02Yqz86iqVrx8gT2NN1cFAbtVQvhVULaMkNvE3qz8A62FMDKaIN
uOJTmn+2FR4coz3eBT1W+pa9SlxS4brCnyOjAWHZ8iCX8ZD/QGYcDDSArJXdNmGl9ZQRAUYBKp7p
XhmouFnL6QDvG63jQ52QmkerS/1NIMfBHVWD2/ebf36iIwyr0hBISrk2w1gtUeBvMYCK8RBPhiFt
7OAWIBOx7/to1wOL5K7hZNkaxz7FpgYDFyf/uhYVnoxbZYxA6ig7xx19zKnQCdYOf8l+MKC/zUjF
RT/xqz+QdPVXAPY+UkBB0Eni9e3ZHOrbdU4kLecu8uume8UUe68uI+PHrkovnyI/2P0vct65d2Ay
57ZAsjkFx0ICREKD9sw8E9aArBjJAPppofUKr3qzoh7Z9a3yzL1VW5TroKB+DtpjlWf4HyEpSFTo
TXf5ZEgK/k7CgJzzh8+5kMUfJjp3JO7fZF7Smf2Kexnia1fuQwglYlO4kqpBc/BUZqcxHBkVNLBf
Gt1+NnPYmUkc03L7YcYHrFB0LP3KEKQums+ZeYjY/aGK0aXZCcQ3EURdAZNpMEizNzoa9T+pf1b+
plebLpE8IupDHS+Re4fqe/70Zb/b/xrvFcqo2rm4Wg7SjpBoLzjcdqYESaoQOnV/9/1cgH8qWTfC
S76+JbN8sQdt0zQ8B6bc5GB49us2WlUtJos/NwizK4Q+burvBxffbex30EcXeJyljjV4FLq3jqIR
0vvinAF6p8C4VE+6ggjwu4uRD0WdbkBWhffc6sQvo/3ooIGzTEXPT/ohEOGamyIjHdiNuF5heGvA
ftH1/2Gyrsi9nZI5EOMYgnG4eEnud72e9GMqfIah6DxVq0goGgNJaOEhN6Pf8LVGuuqJDrgfiy1W
ASQjEYXQD1wXb5+0pDLPg1Ci9kkQnm2tHdHQF2WN/vo5HtKkGdbx5bLDVUXNI1ar/OW5pW0tfCYN
Y65aG4Ci3rx2wlTZ3p2pj+1EnfkhxD0jESWaflOV17PVZYk8tJ/o9dTGSVJX2lfK5Yzri6amPld/
j/SFZB4JcXswxmP+o2jb2askJTViQMoPPZsbOt2gteUUqYf0WG51W8L5o0j9fBG0XBzl77S+066I
S6/d0kK8q6VrjVmUkfabCZEELwz6rJTfp1aiU3fbfVA3sM1Y5+6dpTzqHuK6nega/D6nvPTlgerT
IRb0vT5BZSoHzSKYIOKnxbIMfwQtvXnYROmoVEoAx7B9IF2FOQaYbx0yk7hnOlQYXCI+f4l3HqXx
goxHaDIbkL+NWFrjqMdKluXA6KhaJ1X4WSUjByGSRc9dvXiTxUewhLoy4BP8fznQlSx76NpFqQKw
oP1SYlJKBE2MX7m0/kV/GML/sTYYyXJ6m/poBnxNvr5axNoOX/V65cJCHm6rPIgPVpaSLlYyMtFL
BiSQlcS1p2SU5qDkLfvc+wVq/nBZDAQIrzeXLCaUQfa1KnjndgPgRN3sMfl6FiCt0wRfMRAObCQZ
cTmP29Pai+w1lroMIonyXxnJchdbEmldg9LTT152L149GRQPmXzwAaovleIJ2GTqzjhrqVicNIGq
t6P9/NurQk03oyOirARaLKU6e/iJZnh5J2Fkub60vS5MyxX+jBYIBOpCb6bAGw+czisD98Pg3mRC
fYKRpv8iL4SQLQackFi8mPWEfblbr6hF74uKTraAJ6JVfh3MB+F1Dv5XkKoOKcXq3OE8oGc4O7nv
MHzmkP+lEB77W2kZKaRqzUppRJqqlhsrAPXdj8ammww3EW3nBN/3SO+JV6ANXSNYdkAuUmk7RtT4
sEZkhExrHwbjzwNfWd3saQRu0OaMIdmtL6jJAUfealRozLbDN4xiTJ8TEPCbLZdbsohTzt0DoJ4h
livj7Eupqh8gGU/a6j6P3b9FC6DnUVbYDIDQKhwhzeITNcGeVqhwLZG3hbfU5eYp+1BJCK7m+/rF
Y5wFuczL+d2y2+mHQyQIvo7gf8COiCfUDBy0q8h9PcZ+Y+2NiNpiDv6LAMktO9rdeEI13DnVe8GY
lRwtPPeDG27HNTENqDjScN5jMQuzLIuezJ1QcTv8Ekmthj92D66Uhmp0RY6U1Tdm6xfBQo5SyjOX
vG6RNqJ4wolQjsZRGGz5gUGp0YzG2SO8cLr6ZqNxBEwShHgJYpujmTKATk5+syUYQ8auB7CmH5GX
jVVFA0UDucfmlxgG98LQl3dh8OqAGTnWVcM8xjhdAet8sSO54bAqS1ZULpVRY44pSXBRDPNphIq0
KS45JmXxOJvS8jluCOHoR1857OrhgOnhsYUSrQts4JI2JUBw0qk8kna4VtHoFTL/TEuHeaMFdS+9
gmZQv9ZS64YBzGeMgZh0ebcqPupglRo6WBmgDFNI7DNQedyFlc9wf9ePWI+QklMNAqA/uvrbcTGe
kNXC66zI3XpjNj3YpC0cd9TMvzAC7RbxTejKJnoMkLV44jIdtaQkqD/joe+iK7uThak4W0mhn+aX
53CULX0iLymvqfmBO0bFp/dyMk9rziA+Wmk4ePgen5MMUlMbpFhFRV7vnEBV2vUKS70R9F8cjHAX
h5NuVPecXu781htsrWkHZodIGylGtckW9YEgutCn/QYhYksHSmLAIE9yXtnet09Sh6uXA1VEKHri
hV9xkpkpX0mB9zzaLo6f9HNyzK0QiCVgeVDzfMe1+C5L4YR1tidx/ptdp3HQDAVE8jov5Glc1WTy
AV4QnJZ2YTGKMF4hRmKZaoDUsYaoZkHEeVAFpyjWc3ImzamlPrZJlF/x+Fyj9bqfkxx8KbGPXe4H
mMDMtPKl08Q4uWGLbWlNHGt0BFwNhNLV253DIcNdUkaudePSKISEW0hgjKD2FEwru7jptU8lwsQm
MYbAaA8G9s2mF2bOLUUjmCN1D++t4i2KG7q5d2eQpGwu6LZrPs1BAvD3g81tUPYn6Hplq5xuZuJr
rIM+G8gTaFysBKVkziumw177y3j83nSFeANi/RFWsoyP7mPIjZst9hJBFFuylyYHiDmUwAfSvDAC
rfcUTMKDrmXV+5eiyQvcNK0puapUERXsaU6o2c0bxhzWeed+IaSqHBorpUMXh0L5+JKahAiS78XO
p1EbJHeR6G23cr7iPjc+tmNzlfRDYOn+DewrANBrO+TxORGjpkUgXKHPkUxjSFVleqt2odKjdzTy
f8ygUHLhO4Xi0+0X7WpcR50/1N3/yYlTO/DCjjgPEVh82t8mzksDMPeXdMUZA/Lo+tPBvgYKE3Cc
9mcOLgZMMf7acI4hKVRKaIJIc4pLXYdD88Dn3oopiFT2kyku9RiMrnixR6Fyu3HpKw5L8VEr2FBV
WyklT7B6iSbwzTMx9O1RSnvTJjrQzgcfuuk3ZnElyF7F6p3EeWiHqPdfEnKIlP90gCMJdJtNEvFm
Ua0mTQ2rLBFyGhZar4OTRFVgqywbS8DiidGk/nUDvGfKhptjBQfOnZXT5Yd4ixwtcf5bbYrZZ+Xo
l5AdqwVrLfMKL4C8U9eF5iNAy74vVfmK2jDbTZsPF4rvDTH0p5q8Ub8jK/CGFxK1UiPTLQK9AraH
wOtZfr7SgOZC6N2rU+EuMkLb/UJYLhKYeQ/RbMg9uFWZs3/QWY2gd+r/Qus3NKn594cQqfBj/u6A
/+kQi4VAoDyCI4WaUYYeG1HIgATqWyjmoOpGiIRIpQK/6EmJruLbMOk3Pp0DR7e96hJlN9lKvctH
cximURTwpvfIw9V6/uXV5SQmv2wz6UELlT0CtQrugTIFZJDqYgKGTYmVeDvMRXShXqlWVaI10sEx
ymmTue+/+4sJSWL0d2sgsthsvBoS71knlBMjUr5kN8vcCRmctSlP1gLiQTS7ZhH+1WXrjmtb0fpg
TCxWOkxJAKtKlX3N5q3SDmC06qBC8SsuexiqrGmIde36TGBHXEv3XGAF6UpkpIcnTKivbw5/yWtb
bnggppKa+PKKW1cXnBMV96L88WNXOosBRG8iBhB/RGRiWgGBjip1zwyqr7JCXK0arN5cBLaW97/r
DOjVckLfArc4Ahmrboz0SOBARIGPQ1Hg69UEN5Kr0ORThE+EhW0fW8SPbPYXkw8WLYJD8JyB3fV0
WULHswyjLKjlTK4MHV8PD+Qndf9TDfc7V6ctdd/hwWw7xYgLKh5MRZ6wgXwkv53IDSL5eVxYRF0L
D7gX5lloepR2WEGNYvJydV9X+qAN3UOL/QJZFjR48+RMtiXeGPTrz7gSz0R2x2Dv73rDgdPrhHrt
HggwilrQ+fTgbpMY9rp331TmBas7wET8T8gZ75sqzKJRdFvn01FCTMqD8ZSHilNyaS0rRy+86WxF
wOIXV8UbpwM92tz7hp0KkGxQugwmyQPFd2c6L8DtMAEkCora569bCGag8Ml5SrQWvZq8oyVs2Tmx
IBt1bphiRIh5tpGysq9ENVgC+vEKjTsN4kz79kXJS5ejiPxp4tzyNzPGB+e6xvA5QEEXLcWWriIp
N8z9UBjD9X4q8OlK+BKF7hw9KqTR6L4RvwtjUnchAnuYkxBXFO8JGq/J6vd9rPnGVNLWgNYSCbKg
h2KbHUDEU7ZgcWoEA/T1UpZH1ctLbtnJTrQ68YJ7tTY4p9MOvQNzNqmC5/0oTYEml8jguLCw+jJ2
BqaL3WQMKGggEK6v045urfjcHv91wjnikZQpULb/sD8mitdIBsa5QBlVvgHbx7BM92Lp7jd93PbA
WFA3KB+9gF96ssRedrfdaNWwTB5VUz8eNQ/ixfrujwUXTCodetqci5doHHGsG7bsD5ycBfg6xkmr
wyMGJMwHI/Sask59r5GRN08/D+cPkckMpzLaISi5WglnzxnC8JZO06HEM+zBNEejx50rwwvw8PLt
l8e7ke7/CqzISL2Ojyz6LspkSrCEX7/b4ktT5Y0kQcLUZBZ3sw1BBjaw2qP09PA9etoyAVTq5/0K
+x3rQp85fjUglRanyV2HBVXj7REGh3UIfy+yfSMfFUxEr2bunQj0MlIWsObeec6pdwBRdP/bbtLJ
Owyhyamlnt+qG4RnnLFjeQjKNEtlJTxHp0EnG01XzoTp8czvgjbu80m7/6Jt4F4NeX/W61GL+c7B
2Kd6LcA1YnjFNN2iyLNR+E4TAIKqgOo1Cvr0dH5hkMmzspIZHLgKnSfdwcI1Nw9JKS+FxhvECbfS
wBcnUju7bM98asOVgJKm6S5CbbO1UJAQ4ukXKrKwZ/kDU0IcKUZdi2R3ahV3adVeV40nNevTEPMx
ewWS9gi0KU2d4boYJY7ZFu1insspbeBwMIK/pppYtfbyBHQjPzvrQCCdREW9lqrgD5WfxvQ2eF3G
l4CYzccOqbMXnBqSkHgwzPKiQNB/kAiljSS6vvxcQcnSqfSk2GihqvroBNk91Y/TBipFK5Z1WH7P
Y8f/lKQvptawLsUfGTnF1sFDGVWeXShrjeZ5PmM7Oi7m2n7lY75q98JrWk5YaLoUtcuSVWJmkYGQ
ofc42httG0BQntcsTnWtNd2Zp1eaWNOjemzadBFmS2adLtL0TYzLczeqCW83TMSaFovnWgwRS8xG
2aVZ+rI0wXMFnQbMPnGpMtAbZxWkKr66UODUpjHhl83KKXsIuSUyx3espYFlxaogXnClqEy57eN6
aXuLMRvbntuQ+VbFTOaCQGxFGIXz96qhyBJFy1EQaNkcA3GR+sYjNOk9Xh0RMxs0j1rPoJhWCFb1
N/8QjFj1EwSF8+wy4Ltgbx2+2ORTTu1fL5m/vpQd+ieb43+LTTM20Y1D2P89KMClmU5/AMLlJ2/s
3ObHue5Z/tRqCYUQ3SaXJn8uuEf0UE48U+eeTNkpUCFdqUKcS5c1cj3ML1FgXWLz947s9yF9xvjd
hpcRP9aYgpIZDy0f5jS0XQISGJfZ/x8eCu/6fdb7l3HRuMHm/J8SlQPQtFtPcaOSMGqJxDotrpoI
fPbEQTx9tPPhS+7Ts6GygwBaTAR7I5Y8OD2siJ8vgUSMB5JrAxSAj4Xk7B7c8LLnPYWJVgow/79+
M1xc5/POohVxB89YpekPfoZAD747vixDCjLvwzZE5rFAhHE693Y2naWwqQACXKtGoJigONDo+xxD
Z2wjUnQwpEzyoonlEuhMP7wuoNhNF4Y/PPcv0uhVYQIg5MHEWz+oCmTykPxiOwMfwFOyrHmQP4nk
iY66xVa+yTjrNUpexAnhIdM+ty/UcyE40p5GsvWeAiw353Gzx1dsRu/IS54ROmVhonw7J3XtlJ1F
czq08WG4NIS4h7ymrHi08ZowohPHLQ3D+p8RBhObo/J1JGpMx8ybizYZFH4G86svOfvbVaq054f1
KKGj4XU/vdCvuwXAtVFuW6Z2A/E6w7Rm1TLmKMk048Vz78EyTlVUR+FTlnNkor9hHqwSAK4KdXA5
ZuawdKqCBPKlI9odfoUlzGZeXV9ztiOPUUe9nI4L9NFNS9sZnszoIOu6cYpfVOUiYgbS3/dJZ5St
D2T3FBD5s79LtmXFCm3K0OUpZwegzkF6AVMXRy6CaRGpKrotTXvQM0r4jNP3kZlpoZ46qnRthhqN
Epv+/2aYiI6M1qtqt3C+lSxYYJwvT7lCmhLlFnJLVy5VKj7LmzljbLy/GfrpGP528htzJdZU0GWQ
+MQFJxgCgK69LnhoO7As8I2AcNSi0Q7We3w2pIorxK9ePeZ8Gpiy3Ad+upRnN3KadmUNf/zQVsf8
RaEkueTke+QTajZantpY97K+cWV/ld+pVhXYoa9qEk16pVmv9bsChCUVg+vuDNnZDpzo6+pCsF0U
gHfd3vEVFEoYoT4Jj9D2gTNehYmo+97n9UXx89io5rXG0dNjSnulTFQJUdhTREyhRLDE3Lul4LHw
u+CSAFGanbpCnwT0NuYhMqdkEsTwWVHFxRKORb207ONObeMnv+KRYYoOHZ4u+3DX5FbUEiR9za0b
oYn2NICfQQ5h51VnqJrPBOz8d5H/XiMN30VrNYAyUjG6rCWszA/3R0bxJgk0aYwg9VhmGoPHHG9j
pxdcm/smI51qBIIJmDUmw+xMJvVDiL+hnYiAU8l2O06lFbJLKqPYIcm9yEsDPwNiN6V++pHcsEyj
ozjbYD+yAAKswEEXA1Y6bEDvU4VVa3YaKT8M2ZAVfgSNmt3RUHYaTLaUMfn/bsbZiZFK17YUZV02
/QmmCjnvT5ItSFigsAqHzDzshkTu8DoRe40NBZUWNuq65Xm+bWEikp9wokdVpRirhuVbq9n+eXPZ
Z/VuhBymlHA+xF8s9XnPb3ZGliVrvC4wb7R7qX1s1rdwSpeAVfsD8OiUHSQcd3+cDdA120B9pQti
uxaZfZEMAgIqcWsptVOBtS54IVXxWzdWHZLyOBgLwK3Fl+kRwONW8gJ0Zyk7uEFttokCcvjYWRQc
BwwItQQ3iz5Fuu8VRn18xbLfH7Z6HZoh/e1eaPp6uH1xUxKG20JiqheZ+FtTwuUyWS+/olQ7XiD3
q7wT1o7tWiAmpxdjCQ8jfUkDbp+Y/zy4VqzY02Xn3I0Zx0bZyUudlcz76Wg1UvXA8jNybz8STssb
EnrscC5Ky313PRgCqnHcKZ0Iv9A0c+E9pVE/PN3pns2zLTJ1Hs12+TvcJX614XNcBjvW3YTQ9ZcL
QMoVLiNFw3IRBC3sKtMuIHhz6Tv8bapEmVcIahgwpV/70NoUdXm++DBXkWE25Vrr6+sB0XcM5VNu
zOzsToSsm2kDvCPwXt6QzWoQeDALidZ+MzeTAzCarpJMQTLbtJ1csDbZV7rGB/o6YO5dViCrvvsu
APN4yAx6PG5k53lrozOXYPahNRAcag2JfNvM0at4Lz5JN87nDfAdLUWSFMBORF1cmlidqhXjat+c
X7jzbW4ryO1lFF4kExCSWqrhfPtzXeCTe82XHS1ga64oKhK0CRXMID11CUHpgRRi3BicCS+UKPiG
SCwWJz/DJNPURC20AaZaGmk7dZ+TTKa2gt7JE8W57ZTm8DZzY7ERiZ7Ky5/45if2zzHuD5B4urhy
HZ+XS+9y6Qp6KXBfvbNfED+GrtiAihq6KlaHX4lg2lXN3VLfuywZ2eeYOkpOQZXhSosk3wMJePPg
JX1yp2aBZR+BgJpmBY7EMAWG/y/q+FQnqepU6NblcM0+fsejVDp8xW3MEguRL60COdsFoXOd+0Of
A1uX36wyZshJww2SO20xwy14aE2rK7BqMjZkrTVX6/e5dfELf5DchzxbrSOAz7hnbvYXv0wDioQW
TcDVE8BgMh+zzVzYQxBiN1gmEwSfFHXQtQarwrBgEgerNNjcrncn5+usmMEAM22WE0x5193JRKp0
dal2UFz288gZUdMt7vjhWxd025T+kjU8+CmshMsU5ufVhS0BML8jzopXj5hl8lOuwsLc6hQxUuXw
oxkJVxNDxi0z76JWy7Jn0vQpjU/52Y5XMVN4T23+D4TwhBzjw4ulwScUJkSoCxnf2SKwcKyMAuMC
9QfZ/BoYoxxVE/5w4A1QDmkp/Ltovu7+llZxmjpB+awCZta4MZQB+wyPMl7Qyg4DUdTPcaPu9A4S
vMMHkbGAuxlFeEs6Va4romG5qn/MhhxXo8cMIThyBxPyvx9fBZjA5t6S4yQA1tuCXzS8tzT4tegt
eAlGQqprpMWZkIs4np53UaT+XWaohBMdg2fqo8VCR+H2MTJCmBCt6ecavMutU0GZBQzl+3Pgg/sz
Fzcp/4e7ZjrbZG4/FvaTidruskavELQWPLU6NirnoonMU3XFogO2T8NpI/m+zbrg4TOjOuQtS2lj
5uA43tDTBWhIbnrltCsVJaxTuo6XE8JzzmHNPFUQBzQFzuJzUgtAn3RrDMGRl5vji9NMdmkxiSBU
2qF34cNDCSM336dnLhjB+vOhoeFniVUHU87975Ehi5BLoHPL9m6pm1NCs0EBZKzBrrkIJXkfKtAx
1a5GU1RW8J0mQnuYAZ69Ib8rKBNkg2YjHxkddKBFbggi056eo6GmyZJg67x0wqKC1UlJlf6W9BXQ
DBOwIUzwlR2c0aTm1o72tAbbKF8BtD4t7tzTuuMIvTm4HmiJ/3CPKYRRnBc/r1HeGQV2qTTfA5Wk
NLN0oPMzV9VqErnPzOAvDdp68YY4XaRRXILHEKpufXovqo1mZ3G6olnQWGnZ3cAG+2TwWo4+IpBX
pPgyY+icdFNBnRh7n/ghqsSUDYcx5CDVuazkGk+eDlJQOMshYHfEQf4f31izut81LAkIeC7gr2Bj
2AxUUdXqgWAB1BV0bybO/O600GWzpWQ3SDwb36RveZvqWdCoMynhaNROLaCQv9Hf2IgMh5lGbTCH
TWiQ8k6AmYSBRIlGmZr6iQLfxn+E3nDIEt9Ei78xwRDkTfFLczeyI57ryRJNa35QRpsjRrStpJ2S
NGYpBqtRR0rkHgJWe6pOsxAQ+vW4JfWR+PxZQyxMnBznr+JLPH8NTbhb2hqqkAr97dPtGsTpzotU
YIeWI3DL8SVOyuw1kQdDWZL2gX4TC9aqjQP6wuIy8J3iZig93eXlW75coDOEODTV57MHEcR+HCeZ
htTjB71Wofx0+K5eCoaYORSRdshUPQn3ydt9UQYiG/PGgdzYV7fukkQn8IMTWW+vr5oRp8v9PNbf
OvtCm/qUvCT/XitqOARBLZd0ZsbyBz8M7od9Ye8+9Ylu9AXph1/Id4w/Sr/ErUE0xzeE+tqMXV/X
hF+9mraED3tJywOqWWlucOI+Qnak1eeRlsewcGHDx3uiuQuNKpPF3xh0EfRja2q3dBySCbEL7rd9
6kAb7zTkaCh4QFBYx5QNHCsfIMo2+DXBC65aur/vfM2fCq0MrMAf41aKX+BaZoBKjZgn1/CAPTzz
6fSnbC4e4Mw+K3JBccx+C+RRKZfM6qGTihpi7sitGkU99orDKzE+Gv8ObyyLDwLFcE5pz+/Ksn7F
puH40SyDkCXUSZ1rjj6yFw4gUdGPis84ehMb9y9Mmn371Ez0g1eszqBctEdpUC2caUWN92MZ0qc2
nGPej9fFRf1NQtaEg2deKit6tfy1zxBz6YGTB2XlWPsjPNy3XguCSxzuMOQNES7bVwuTGtZ1AE+2
GntCgza8Q+HR6RVFvbfqMhciU/KC85R9j0r23ch/u597pkmhUqKI8THIotNTgmjMkJUZ39Ul9vbo
ULrl2m6jJUS7c9Df8YCrTZbnmRY/Da/OgS0zP+7CzZWTtdR/mxd3uOM3wyshrZAo8EyiXn4u7oeG
l8OqexpZh2kHX9atSkS7/gmEHj1wTTc2nAr3htZ9zP8rLcv/kXFdk9rPDedtB+EtQovuK3ga2dQX
e2NUYSp25Mg/JMZiokoS7WKUG2fPu0FN4bNAZHTvVAP0kBWR9UCTipSc6PJgeT2naxAdRG/v6DnV
ocVKvkqW5YbhM23dT0it64cjHpX7ysEcysZlKvmYMiVV9108O1jDig4w5NuD8KtM15WynTxQyYyO
AtDHsAdbkZG4JQ9yx49louRgHBkYKzwXa3wKSTkJZDQZQ4ysI3uygbqaZldpmEXv6X9vTpIlJNyq
meIujKGs4As2en80i7UGWaBoFhXHJbPGVWcMkIWrwaBVyJeoCP0g6A6JvapfiSNQxCBsfoJW6ZGb
O6ZS3fGreBTB8Oz4sO4n7SzrIF4eJPIW4nw95yLvG7RrvV0TrvhWAaY8vJzFVbRH1mMiDVgAQJ7B
ASb2JChxYLTgEjii3G4sW25jl3LXFHHMOKvu8inpLaxLyZJDYcZEXG7Ww+mR1QLtvnCWgyntVA+M
AcW5/pL061K31cXjXYTqya3bt3d0Xp0CLG3MdkyChmX+IYge/rjg+h16llXTa4Ru+yb9gNg4QFD3
q5bSdfQdDxPGVwBIymTzmrO70J4i1ssaU9W63UYsD+YrYb7kXKO67/FgtosZHTg4mO81bLVMdKL0
xuptNjLWJDKEbo91QNdd+MxOMQHf904Ue2TbmiA9BPWwPZHUOFwtBu39H/TP2Gpeo3S2BRaq/wtA
+G2PFJsK0tgxDekBiqRLp1r6YoFNSuM1Z3QbX7JOvjOlmojfCP9qCp9/UUc9eNXnxAvgQpPNOZGc
V4bnHXW3rgGlQyCnQDR7DnJlMRTxbX8+hCA/6Hfbg7JLorQovKrCONRw+akE51su979mkbgQp5+1
S7RskcnJj4W5giHDZCukPUYtOBo47ItJpCx/KNtKuhLJkGdloEAVci1DBAzyi4GfT1Iar5mnhd3w
CpCJnD3Wd6QWmADCIqH1S2q6lhH6jzvO/6c6xxr/TaFvmNRR4d5/7vWt21ZNFZJgiIiWT3MDN4NY
IDE664S2A0+duK/ELjEMS3PzpAwAR8V5F9mFki0puVs/DgewqRPPTZPiGaptT9nuxWrQaRjhTNcW
mpBtssZzRt/jheLZ1wFdoYjfLuwi6FSPOnYmcsTjN7ApkMNv1ZezsTlAXVoSJIV99aa9DIv7OPZv
s6eR9mkGevnPdi18IhmJ4Rr5xu0/qYQc767BQh/lbSbIa/KUB33Z8rWrG4TkDlzbBXb4wm0gKNzh
BXpyPKQQp2OVSfzuo/njaDmWcjkRK6chIBZTuG8uwvPXyTtOcyx1XCNH33c9/IZgOTioXgyKfeEp
KEq6ax0XmGWKPPZWl8xsL0WLtXwtr27tllHZI/YhelvbStbSSH2P7XX569VGfg37yVsr2+JxjTpp
WFzMs5W3qfdBNI+N+VgGtzIDNLOrFTOYm9Ay6YgqnfOo7llsg3dCNWqRrH1UvyLjVTsK0XvYpXx8
5iVZqwqvoFuy2G94ShV6a3JPCUtSu4o6pntNIpmrAN+uWyt9pGO8iewJB9mzGEO3u+JjxdAjvB3k
plszNwlamaFQqS440TPdlGS+AK3X/Gi0eCphm4sBbgul2Sh/mEjwBz2P2SsJd4dE4PEy/7SJ2o8m
lIUKrs+oAd+Qk9c3wOGDYej0gpitEajyhxlfgXqzU0SAeTcBMvBCcB/+hQPJwh3LfkquPH3JK6/l
ydBrlYtn1EqIamlL2igE2KTDgxJ5zpsN+r1pUna7zPHgZjLG1423hOp8qE0PvgCNEqxLNn22npsJ
nLLtDGK2jKLBicke7BezjPDmW1jXGXILz2aPsV1NtEPHsZg02zMiiEuxuho4xwXommbghOdy9nfk
7VMXGpsNBM8y77Uzs0gIPEvY1HFKMCC1rV8XFnhx9FekK4mCvLnouijIrhfk2KomOUL3MgxvSGa3
VEafG0JQEDOFcteZoBjFr4so9+X9MGiqSPdkm+R7pXchtifR4XxqHghT8qddcJxlPAsJ4v3vifb3
9eB7d4g1SjrpNik0iktDbP4faHnD3Q9ittTnNG3Nlq9KsqeyoTFFnP6xfRU93j3CMlS0Y/HMgFFX
vg+aOPMu1l6zfqEMHvRMbPaLZaeUo4MkfhlIgtAwXXn0H792JHnfb0lSCX7HyYaYd0nNj9pOjKUz
BPwzRPEM3ZNkr7/1X3kjAO+HKBLb2XxOf2IdJPawExU7XRc4HJEHUdMDWv4bHjl22yIfbP2rw4Vq
ILcj0TqsN8/sRjQ9hb8MT9+GWmjEQ6/qPLvGHAgJOyjFYPG5I5gq5nKppYz6B+2EkT5sVcqtL578
dPjCx9fzPyVht1X//MFtO2xmmR+yOuQJTTQY0zvXDEUW4E3rOk2ysaSEHa4EhX7FavDOWI/RJHN0
x5DMS6oFWXTHZNRK3moniAbdps9TowJD4pJ0pNdPex9hDBcEzvzIeOvhaBHv1b3t4LAbOl4aayL2
fhzysrQ0UgZx5zo/RHQ6YRR6gB+o9KnKTFG8nt+eFH13kW6IrViVudqBiMddCzbxEKTXpB6L5DdG
/FFTcAscPmCoUCIlFoGLKSVSrc5OUThiDfDk4Tk4hGhzeHZWPR9VF0qz0G4GgnPAiRZyer8hom0u
PGrnHjs7QEkIw9+6rfyA8B8VrVgrHV9mRzcXYNHr67cF3G5qOv5G3AkpYTPilTYLm9xY17m08d1j
9WFPv1mxV2PiVXH0ND3WbklqlUqKkIRduoCBadSRQVfNsn3l/IzdEBr8aIkIVgwtu5HNY8u2q1RL
Pumh8P86vDl0HhiiSwRmtaCwQWUw18V/V4tYQmASeEqkOYwIIPSIKlQR523oAfigjMO44EYa4OBq
NPU9nlnzLZmd4bahnKd2DfC4ZDReTQwTkgQ2/0hTI3r+XRT8rGqGZoNKW1//cxPieqmF0Uzvh/K3
45Y0fmHfOw4Uhma1FaODmBhZNFrSfLrOSuq+UOiYnsFMEr9ng/0fdfJqLZ70Mc6wnydlvyXWpiij
A8j81BWy32tmC67sbnWFiaDtNI7yiV9o8KRW/oX3LGiDEiGMHV2uroPWxLJOrVJXdgR8XHVRmjLx
oCCCNsGePSj9lxW+XxB6Px0VGLWgDu+PY4OkzNFguItBZcpYNP8cVkVgohM/b7/5hhMEzDI13m5P
mYFjKIaRNRZchP/zZImJ/UPsLyJBK9HxYVA1OQg39HmJjqM7w7oIQ8XMrgi4wUNCYvTk25CQChJ1
RPkQZB0eCIaOOC0N4rlI2ftN31fHsjMxRs82eFTA/hOdf5YhRmdkaCM7cMJ2Q/JEawmScPB/rdf0
p7IeXJ9iHuGkiFtkzwxI9EZy07rqe1CgjttjjAqUiBw8+Jd/g7HfHO7JWXBjzSY6DALxO7e3WuFc
CTdLaY66Mbf0mibwXXTi3ZUGJcfdCmoRVIIFa7GWqvCP9oUyNglSD1hH+l2Y7dZLqwRbQq0vYDSf
3JlFI8P7G+bPDqN3mZf5uksYht6nSyyvkJBDAAHbtz84YMam9NAjG6ND/F2z4G/H9lDQOrQSdvej
JCibzmfeXxAY6kX9GYxCczkZJG7/x3UGXXkXec2Z3KMQ0Br9xNv818LYzIr3ov/wTqt1Bjt43GlB
lnJCd8b2CotWpgzj1xifm6qwYq+g4gMZkJRkhAzAhJSGa6UwvRt4uP61PE47dA8uEml7vjpRq/yf
1AHzFarGrWTu1hacW3tk+Xi7VC7U6KuyLOSb9ag6OF0J2mtno/AFM6Myxna57p2K1Gyoe4SAFW2o
Beh+afTeiHhLNmGDDz+P9xbrdMKPRyyBp4PARY0NGT21T0pUFAuv8TBdnmoiQlT9YmNX73QYdMVl
JsXqZZi7BHoqaYUrRHKrNysx76SwlXb5cyC+2RI5iViDUp37NnGUXJOz6AFGl05eP4zCQQihGD9u
LEh4IERw2oGxyCaTHixYKJB2trq+QkzdFCgqGlK9OZGv4lfR8nYge6blNw5zHfy8H+cd+3esUb0i
kGu0tmZYhcCczr6ibFk8uMsvL5z6Bf2xxxoninbl2I8IefaFlaQ9UM+iw3B1obTlPjjB/cJamOdb
3btuTvqiBDaXDt80c7nZdoSlt+WqR6UWtr33EbgAsngG5sPKA3XGcqtHonqc6T3A5hLKAIsmq01I
4EaSf6ct8py0gfyXDF1JCLbwfIYFIyI3leobb5IiE9xKFFPFtWPbsw3GljXUpPtbywaltyGhXpMc
qnM6oGJzkCv4Sore6PXPIxSNninqHeh1Al6bYowOjJGjdQVct0ZdgE8BgGwYiXbA17HtbpdMhwk4
LHzUvLJoh6Lh+TgiOLozw3MrxFJq7LIbrSVzMGdxOrC+YhFp0vYBvnFCzOcAgCeU2FSREc5T/LGR
gsPzjf93PawGrQCAHKeSMgJgvHTrwG+Cp4fq8wE5d8cLWHq7ZN/VOKFKtuw4CKq4xkddVde9ZLUC
QI+/Of67XQcj3yqlE4HTayt1lA8TL2TgNENYPtJG6byhl/b45mZ5ZoaxEoqZZswhLNNc+/zRaMFt
3wp+EFoYJJ74vJnpRJM/GLQioIh5b99FSWyGo604WkltFnryrUPwGMgHvJCcSau7tia+j9R1yKm6
+0fnVlAa/jpj6xkDaF41JM5is9S8qq7gw24kDVq+2Mw5tXvC1DFS4xMHvJvjiCpvKGTfLsA+ShX6
GhpYZoLaqYi4GnJnYW/XCmjIu8D+8gv30KtrNoq2gmdqKKpF5IltgkZf8G2WlcVDwgPkjFydcyOI
o0S86VL+OnOfWPeeQR3FTYhCn87RrQY01RUTBW9hwyRZjsSWRWbG9Sj/zzkW9jarXLIq/yGxs+6J
QD+uOjPFkIXvfl/ffSrR2K0Is3siAkcsM+8iHO776Z+LbjLjjYpFDmeaPKRJawkZLRP7On41ScBh
Bxf80l1qrPhlSHW6uJ/N/jy5/BZ3qUsAg5CrTvHL3tMsByvtoYvbfjj9zSgdU0mBOI0sKMASqqyd
YdcBZJ/+qf3yA9JZv2WAfOJoVvmEvSGAZ17vvzq//6aVb3pphKtDJkTSqHYehEdNsH5EK7Ia4W/L
d8dbm00o9Gw10cT+BUNan4XgxmQf4vtR3dvvt7oQpXvvGh+jt/Jm0z8pmSRAjFKEY94nFYoZhrpP
IPrMTPMYRSKF4lghN+xLkEB6FyvFev/WGkoQmxNA9no38UbMlcL1E9u3ddXBp+FOOAAOWmy+Q3cO
JQ8OlOt59oACRtg+zyn4kAWxu+ksPYbAzqtKMKudVVxpfi84YQoFStW3y+644h0/N4ApdOTv60Ze
4CfzEPNcUhJpWv1U4yl9w+EPO3n6iG2q/sW2yOqWjuxxjvXcEGjw8VMPhMwxalzAVcXoWSm9hDIh
rI3xUb6SiqqGiLmI1JKDGar+bS29vBsQSxD10hI+UV0pGggDpx+wQ7ar4C6X3+BZI1pyjKMSOnmK
CEXsS829sgBfsw5EQFDBeP9Kgc6c0Q1P3VWgTUqZNW7o7bhOa2xDQa3fZkrHQVBVs+6OtuxjHrwV
mNIp104mtusbO2gBC3bcfmK3SM8Ef5RV24Qj/5MZ2Ea9W+yO/4Ng9SALV3zKPWn+/njdt7pRG00v
78S4Zmr0S/pdo8SpEkfF9BtspBQJrlrFksLC72jsmw76dPJYHBw6JsXJh+6v932hc4iIiXizw5VK
uX8gYLoRWCJrPSqnIkoIn7htbwG9VbdjHvGgkbmmQvh9XNJRCzO99E2v5J/Fj1My/wyiSCNFl/VD
6jF4Edtp5PEwr+3R2SV4YHYW7MO5p1Yih7tGiFoRc1OPdeQnKN0wj5iaSqHiMlBnC/LOtBUK2BL6
uvuA3/3T/rzDkDmvPu2b+M6VRXEXF6kdd9PZNdty/SEZbF6wk7TOyMh6ho77RJcgoNSjsF2CEuKs
SA0PV4xSiErFbCZN+JzAxEMz0I1E9GqVOVGvTbyHguwH2UnN27RdOOdXJ/KDoGyDcAFD5stp7PWH
5OXXzYKHwbjViWilZyBjPKJJHzWBCUfct8oT8q2TGNnSslMkYG2n9LBbuP1K6qA1Nt2bOtiHIc9R
GrNLjC2veeXC34UqZ95AUkIxaOK1Gej+HkJHlAXc/mpQEB5N248blOorTXTfrlMjoTX1Zm/WMHdp
+f/URjZNzurgYGEnVHxXBaBCVoPvMLEy/ExO+Jh8qmoX636fTnoQ+VMWupI5Ms3ynsB+VNyE5w4t
UDB3zvZtzpyhWRZSl8nCJE3i0uRsPKHO9LQ35olMrLCWArWA9lCvT6GQrYp/fmNsOh9HWJEJZvqg
pHEkpu0j3qFhv2WjQ4aEvKMyFR+YYfgNkuOoUoKpmd96FjL319nQ1DXAIcINMQtkjg2V9Oh2DvsS
sd3MAWVjjGU0ifKFmdGGV84C0LWVNw8dXLLt82aSkCrs7N5N52EwOs71/V+emj5k+O8uABp25D9L
AGsaXQaGdp3qs3js6BxiJhKDBZe1cTr+/DiLrhDayLwXRPeuZ61wkVQZTd/F4Ejiy8xyv0NTT8HR
1MSp86dRdkI8Jlx1yfkVo+kp+13FKf9IA8Nv2eFj6cG6/wnvytlAGGSgEZ+/E+Yq/mDS5KQhIbZQ
6hl+zgbkTnnbcm3hnnaNv0vFqYWRcYFREJdK2ry2frxbBykT7keWboM3m0CTgVAtnc8ZogGuV87Q
DNMMpaUV/JU5woYt9/s/DMCD6CXjTAgWlijQqN7q24j0Lu2j5eD1O7zCFHgNAkJu8Wiewuw3Arvl
DQ5eJP5JDmKA0gRYX1x66mlHcGAn1w+ZDgJEYvGKnAZjgeF+ursVVP0a4sCr0x2SlOoudYgQTJqP
x4BO84aa1Pfe6uWbR5TbyV8cY9F3o+QyqQBcfEKOjqyKARl4co7gotUk1mzZP6xVdsGrdf72RP3z
5ion+IyJaF2R3mY1S7Znz3iJUQmxPRU8iz4DaYdiOTx6EXpXUOeqJbeeMZZY6e4rywpBiUWwTEIx
uwPZX7cPVXAQZf67tgX/H/FLC5FfW+vHI6MWAGVTGOrnaeNnv8tqwTlWOcKXEmewBdJJJv/tRySs
lYho9+sHcBtaiszHp4qggiZ9Qdl3esnMJTaSO+n7jVdb0SUYYCsre/ktfHt3/3hS872jh4V94hVn
39xyaqjyEfQQECFIOk56pRZpxFjs7Jluxn+a0nE8FHMfVCvZLN4HCbVfhWY+OgOi3t/OFghm/j4M
X2Ncvj/O2YOd4XbcBRNIT6KhSadTmvGOsKJZJm5wjYUTiYKYU9x+TnSeUThVhv9VaCM41q4eSJq6
/tM9fAuSYXWyLxshr51/Hk6FriVK3DV1/QU2C/8i/7IY/UZT4qniZoH+bzMsMYRJfPTKXOAzAO4r
kWuhjxzc2jif06TpsV3rvpgJUR4O9kDE/ZFWcbSGFjswWdoTmKHjJdUjymqygrnGaR0NZ8rBDHNv
EsefIu4hB6HU/Z9XoGHxLisXupUjKrWkNUFkUkJRJIzxSINIFxl0zt2wUlran/ZdbmS8Mz2C7ED8
i6h53vT1rCVwfNf/T4e/6IOs8iKqzSV8jGCdIkIKxzBc4a0oTUreFpkyCe19AAjfGUQJ4ekP/1u0
wt15pGhTNZXLTdvXhhBuaUrz5IdtZp1aLhKjXgCPqH29F8/PrIYNcVBLiJc68AZaiI4FAIHjoP8+
cEb51FnIW0/BmZtqOdnYBWRwU6xeTMH+gfsn9EdeEjWFemtsNZc4Omr+BrqNEMS/C/ebDvp1uDsU
F3x1ddMqwf57+NwMYYgAEeRnjDJ/fpGS5stC1u/7UEjwPXhn4KXUm81saTiR6rUC4KDmoCmSH0CQ
V+jxGgzPukWxN/SlIdafIbIHAwm/To2tEJGS2zEulzDscF/6RuTsUzl9T2YojxhX02dBhzixjNFi
peHEYYyOkQcuZegWzj6bVuP0C70BPcaYM0er6Jo9FHS4egEWmzoRX64DH7yaAsSAD+P9HD8nMVBJ
1Io+FimAmnebfZ1ZDIwloz3Dzv3e5aEztFQWBxiYKJRLq4d3tr6Eioe/J/XZy4b0TNO0Bm+gkrf2
Cn6MadKRgJ2ezTKF4RV94LTdH/BEloKbCBUUrx8CQp02l2YlvRQZlQLAnkhs9IlkOX2vzHmUE2Ob
rMcWoVXqiVz55RM/golLPbsTcg2Ny5HEy/OQeDzeTHI4UgDhijn897RTDvB0hLrQkHc/+N5IMD+h
SgoHFewKV4/vSuiOFLgHi707pCQHcmtdDz4RTkA4FHbipk+fpQzjzDCtpzLzoJE5EEJo3FuGAD0l
z+iZX4SbXcKcA9piSIRc5waOybNyl9tGuHeDri/vW3b0FeuK3nT8k3RXOehPaaCblbjXInR0/68o
dyoka7l/+wmFxkFn8n7ozazUt5YBPRAOaY+ar7dtvCShnoQampcZF2XQcVm9yGY6KnNS5esQXqZI
dRXTcGcwV5MULS1lrpVWwdtLzA7K7OVTLg76viUHmiPZAvIAZldw3duh83UPXEeSYphks+/YvlAL
SJT8DbiN6XSd/66em2QgqY0o+96DmOkZDJNMC/6goce3PO/YYuKNFKzanP3RrRLMAux+hJyDSRtu
pKvHpdEFPiZKgX4rxErSN8Aem7wtIPqZAby83z7fG0VkQJ6S3SW+k+NtUQnRjeBZfk/HKzwj4KQC
IBwyFzG42XSUB7GEO0b4c+seLd0BFeyjHZguOdKibYq5BfmqeK64OZVq4jgCnPpdCNltVXvDgOq6
gnSIMUkJmx+fFcLOHSJ6tY9qJYk16KX3X071v58qNw1C2LZI95PGEmxzC4ccEvYDwMkPwPCVXAIU
wbkJGAMnt1Ep3/3XZJhOHSz31zNxVOP1PAUf9qmDcP5FaZlsAMLSK9LRkCRuxH359TGBKc+1STw1
F4twHwiGCEvjKDlb1zaw740OvdKe2fiVba8LZiiFLgMQDML6i5ESU0VpUD7slw4hZsibW7PrJwMn
cGIjvajyQ4AhewcHwD0rNpt3XTlJknG2qaCw2q1kD6UkNwSF9DMtd6W469bNbIaJRd42VnvFKPLF
EOOFg8P1eC8bBa9dBUwXLxvpHUbIFJ5HJeeQPu3F/BRZx3Hs26LOdLFOjpb5t37Fjy3LjHLrEFzX
JTR5fZ5luueWtki/0HuQNMfwUrlUJWNStHYhPu/Vmd88FfNcDd/AiZp3efQ6ESmSSXIeGWmmRdVL
/v46Ohud/nys10SMqRYi/dvCA8Q4C7EN9DohDcTVn9eddLPvgIpNId1gyD1Md8wQaZdcXva8oWYt
isBjt8Hu+dFoCdX4qJY176EayyzN1KJeaWrr48ev9N2gdnNCRStct6Jk62kGW96gWnLas+6VcHPP
XdeBVTSK6pQBDnT8OsphyizBLW2bTHqSzQ8Tfk4RvT3/f4lZpVvbMQ3/yZ0YOIOIluIKbD3VwYXA
bowtVOv4/gYyqG0vqh7qPTm8BxJHYeF0K9EElWugh3uyLFsXX3qaWrgvheMtzPLN57s/fncLeH7C
XdI0uascSiUfSoNWzmpnYyK7OCw04sqD2iKFtBxqGDYUj/DMLH9MF0MKE4mu7FzpH9NX6+bgTLhR
LznPfDyl39YaiWYhN7djrsoZSSyBdG6EjMpfKrASUrfe7iOgh3/aZCGHH6iA7AOCzEl4GRsGvv8X
ze/KoAoA6W4JVVQoqEmeqAdUGc5xt57WkrjvbMCAY+e8pMIPgz+fJqkxehT2X8+UlF/C/DWd8OgP
kBab4eAHYJbAtvlnPtRtjZFuNmhw9pFmuHJRzkyAIorIPm0X3rcj+X7ythjzB2VcqxnqDCyAY+UE
hKw7dwbsZmkBvBFT4oExKIO9U1OmwV9Ae+XEYabbfou/5pky7hG3sTusgptppbdXeJQ/HRN0UP0t
DLziNeUdXQH+dWjOqgj2h00qhrAEJ0/6pLtZOnBFMstdMBj4B51e5V4ma+yT1pZl9fNQPbPEyL+G
//BYB9/7tpZJXzkwQ6juqCySx16EyA5JSI9AFOM37I8QYQ2KkhzI1DN2RO2rDKc9obi7D+SgAR91
ZxfOjZ1KkzKSiwOUdm2nMsNywNqg9TI3VYuO9ZmteO7N15MMp7y2ssjifq/W2kgVQnO1cwBS+lXT
WIkiJj9u+wi/1vKaATjlgRFnYg4/+wne9+EUKwC/r7JpvOnQFf4DGScP99vG+Hb+if1496gy7Myg
6JBnF1YpyME1k561N6hzfVPiVrl765T1AERU/sSXcXzbalQGq4dItAvjWXj97v+wkPSQmmcCn55V
D7+CJGhOlkBTs29s1/kKtJuYHjKk6mY+ldM2kAxSQcAV1PmnWqZ2d982a1W2BExlkFGg2IhV+5E7
4tw3etnABA5/8lsZwY6wmtK4POA6Gle3LKyGguJf0M0jf6/vwdLw8ei2XGWSVRhauwuGw4ersZnb
fkL7LWvNgkZNlLAK450li3iaea5pE93Ut4nURjTcHvEuJJgTjGkvZJD4Nkdo5S6TqGDyoiPwntOn
EdSguQGzaM60JVzkkOHRLPAjT0gj37RMVbQvjQa5OQXaN1Li4W35nUh4Ne1mnzqoTTH5Sk5TkCY5
atZ2Gg7zFestm8V+Ovkly4L877fEPeIVkHZKPaSZ+UY9qLzSVSzDtL/w5ej53M1kOHq14oS9lNwg
4B3Mu7aaTLliReLQT/JaQQKwGPuf9Ekj/LYJNTCgLs5z6fYR0Ply1K5FaAWVBcRxHjsX7f09MXR8
DQAasDA8sXVwIQDh37Vh0f5cbPOobhc1bAQKyWlHp38puM/UgSXRhbN9IAdTSd5I8AVOPCHlCHHg
uXltzDyvvbXb/nQfY7NTPjGyDcdD/zHgHLJQilt2sHqBbj7f4f1lDIf26YYv8tEv9wApmr5cNHQj
hGegC/ArV9qAelJn1Vq3ZVAGYL3FEvLNeXRkNYdVx+tSrnmGjdh/uIF6TOkrK6opH5rgfaZ0xOWX
K/XE1kkF4xoDKYSvVVHsVt2L8nTtczeMpUGgtZSjw32OQGTY3+TOTxspmGh1tRVimDj5+bXzu48H
stmP+d+13E/vrt5MuI3lEFa7hHxTu+d4cRY0Hl52BEaDqAn9Nt9Ac3v6knMM43X26UuPTH83DLG1
zacI4hyyJtWRHCtfOQQkXc34InvXfOxrHGzdrFZ+uXjMOOxyfAk2q8KajHy0idEMQRlCxjXEnV9X
fs3ZOMx2kGcnnnUrGIOMAc3JyVUVpfaNDEFzfxLhXv3oUeYqOZujCOHQjZ6p24IpZQgWAUJRenCJ
CtLGc7M652y6wibSc5SLxYeg1/2aFa3kPkzocwB5jODiPojWL/jTYkOLaRLOzyrn76KL2q1BhsUT
Eqka8Ylbf10LfwWvDdFGwpbXmw6n2/6yOQGkZ9Ysouebdh1ikFwedPg/QEk63rWRbvfnt5G+u0o0
9ee+NkSjSWzsQP+7Zu6HTsp2cIQFc3pTCLKk5HCCeVmQEx8qLLc8f9F7gTXEjgl1SsuHqpLVo78C
eDcGhJZEVifQbN0qyVBLqAPTvYJNmmc/DyOEnxLFBNqBUsdInzcqIrEyBgddExR7yeVZwCikGb+c
pDgPB4DY4twd+M1mSsKRDBNyMtHCPxTXYsaLF7uIajV065vRCpJnl7g70ZxF6vWtkg6uSJHl5hAv
7uPCCZvhl17zmn8tgHNqov6YYE/87eLOSGQvEdu5PqbpK0p990El6FucWERGmuMUS1l9Nq0LZFuh
mi1hOCamDeVMQOUXpPzulY7G7mVvMZjYHXHvxORYLaTn3vV9axtw8u3XNOu5sbRrdrIRh8kMn6m0
rMxX1C0PqH8dtzb6fw4nL2CJqKc8EVvlRDZwamCGk1cpccc/rV6pq/LLYnE87/aJD/5Of+FhFOr+
XWpKnBdoMBxcAZLxnLGr0Mnazwbsudm92k+Jhg4PXuL8IclS8mGZ44YZo0eCVsRvUI8m7XcQHWNn
PP9wSQTyFz7qoCeHpxxyk2cmRzxgFopAiUGY3q3OAxZyY2/MbTBwrMKONCtZ2v9hBMfg40oUYyRq
NdPfF19NXSA6L4/PnfjmwIav0O9KbZDyU8DLeddoE/+kD25H/l0+93PLRFwGA/A3GBkRBdLrEeri
QBfUVUu0X2UnPoaGy1NOTBA+Heu3Cx8Dk6z9O/ktkIQ+uqtLgT3+qOwy4Q+7+Q9AbRy6w76dc7X8
rnXxxrZQr6kPRLwiwyBdIgD9SU/Rde6Y0PcM5cPr4+1u+OvnXtpZENKUDgvruuaq3OtNMnGtZcEW
1MTuordwhULCZ//gbCloR6wuOINwLEzHNTSdKmlAc7C296hITTvtIt+otKWv6oIaIYzHBDqF6mnH
yR7Zxr/ZMbj2F0bwV2AKK9Z2LONY61khsMkg/WFgB7XVKk0ZAVqKXxnOow3mBtyqIelgHO8vj/sL
oWDouHyB7WXc3Mb9nkBPsehd9GYaG7Auyzbb8Mx6R2JKVczPdKlL9zoS7rgHW3/NdF9c+Oh3BoFO
f2nTzWOM6ipOQc98p1kLLV+0GHs6htwfu4hjRW001B8TmXvpGIjHKIi0vJ5FM5EECLbjnykd9dL5
LFRSb79+Qk1wYa1mYzQt1k+NXctYiHLGgY/lFLPjRyqMHuIc0wJosKXqpD3fwVvb1UMWRmlB4XpR
9ThhJZPV7Lo/v395CMjL5hwV96ezPQWFnvl9GsNEELDanCPLfutKGOqdY6wYniiLTJuyXuOXd9yt
TyQWYL+RmhLib93uraru2JH2MFWTAggpNNmkg3eHO2AFY5n9btrD6x9aXU6MFMa2Sm0laSNZmthd
K78JSkPSwKU7YgzFPj+5xATBuueDS7jGcC2L4yU9UEbUYpWk0xgLdtvpODxRd5OCdZ5Wp7VJ0Et0
wB3TEUjohYlig7TsHH56DFv7VP4ojUfSfgxG/WMMXuKYQL0iHVFmzbjltww02TcYuikQnQDVbG/y
kOow53c3UgeDL8lK4x95RGhWuVToZOZeluuFqs+y6ZMEZG9tERo0aLYuAb2erz2qifxsuk6mzkTc
226IL84fJ7IGNGVT3gLDRi7wU1Bqmjc7k0RfMRStJsQP4y65kvjo+lac/CoPpmcjeMa02W6qxoQa
A3sqaExsyvboH+j4Ob5Vs3+H5KXAyy7AyFVYXSQkBGT9XmL+LdIZP//QZASmwLtCUZ1jXu5Ye4KJ
iRm3GcmMKfnYLI8SzjKlaBHTkqN6q/fASqssvsOSOTYhpNvkgbmySqsM++l/fpdzC4zRRl40KL3X
C8R5xa4hlEds88E+TgUxIn9WPbaG6BxL2061LmVKhnGJZD5I3eCbq2yoruMowQys5Qva2oJfnrcx
VSJuHnc2yzO0J+2djyf+mm44SDsoWXxX3/zgRQ9Wj928KtMY+qFZCP8AcomyDZT0V0HJEbqueLDE
MFsQDAJb5YOpawiSm7oUnEyaL1X36HuhoO+7Gmy5OzjUyXDIWM2V4XrGD86iME+SjNqiob23usHZ
y/8drd1CWI3wmpVFuEwEc+nEIJ1w+pCMhHC5UwJQ2vEF3UW6GjODEdPhcbYieFb7VYKL941qzYAO
BZiWCE3jEAMyLizFvhx5XAnJ7Dv0m3RfXFGPU/ocoBJpVhvEOx4LLnrKJ5KPGTJa7v+x7Q3i8WiR
+SdusmJiqGVrU30wb6dF6xQxXsYdnkwwrWhUMq7rjzcvJd7vZuZvMEigO/6STg9bfhWxn2F71O6o
6ni79ZPhnqwbp7IqDf+sxBBVgqzoMyB29Tup5kHuC+CA9+QDQl21yBLGe/d2ThzvWKTA+7BJoriF
2eDszSrq4/MbHGip4YTqjsJDwZ1jTywr4pYf3BqBIJV/tLH0abw5kqHZZcHODVjb5D/0bfV3QMAl
odRyxxU8tD3UNHX3PrWe6pcW0O5kVr4jW82RSkeR207XW4pNiZKUrreqY3Na02fLlKMYb7SrcF1B
BVVWoun191nPARAbgv8sSERzZ52+6RV4P3S7N7LabnAwRNcYm0dDwMy/7Pt/IxWnwWdOgn9yWADo
V3UkihYzr6Evi6xhiY3DvUxGlth3Ik8rQjJeNLFzLAUiDeJYP9Jy542Y75zq4V9kGxqm6cmEr0j3
ChBo+YRdyBSEN3OiCCdrDzePNZM1PxRJLNuuKThP0HoHoA07OrHL7Chkf81Nnpjuj+3SW/jh2mc2
VK9j/VNnh2As3/4EgIG4v1i7JekXQogtIwb9lJ7gIEPyXzCxLLBhAgwVHYRxccP4DcJ8bLF0PAaW
WI7zCllMnOmZKYoTS47gqVvFVnilR0poP+80RG3/0xNIzrDqilsAH/IDbP6VDcfWTYrGbQBprKPr
B+rgXPvN2tu81/qJVOLQPV6hWBL2alAbd1BsFQG4Ss6sLj7LeVhKG0uHECUBDPSyOaBL3eP2X/fD
XoosGlOfHGvkQ/HJtKJUQsdubAm4L4kqHXTFG9V6VRQgHQitu2sgl0oRPBFvxgxDNk8mrbyOQbpX
/XicRiArLmZdEv0g6vJMFI+fYcUOgAH7XxSr/1kHJld41qaCiRFCOCVFa2+YlHBMYfMDDpm04fgX
TYntowkXFFPvbZSa9E/BATIT4gDhmQSZ4YxAACucusPjVZ3swB2R8V4kHkio0ptB6GFhZIUHPo+r
OOfDSk0IHvDq73+lg8jtM8VyJ+rjpjX//RG1c1L2T4wS460TRIrBBDeGHI4MvTYGnBNtncQyYfHd
1Xv5EA5zYqo7LBYAgwarA0SgLAP3IsGjoXRJqea3Irs+xRWmd2zbPUe6KgASQz1eQ5qOBBZjIxM+
OJq1TPG7al44FUcP8qCnHipv9IWKOlLnX5yZeo7bFTfIPm/popU+hYUGeDqOr0BPd4TgvCiz1xhI
h/pie65zSCYSqWwuHpidqpy2dB60Cj9OCLXWeImOdXRKgKk9JiSajaX7f0EvazM27hesPq1v6kQK
vC7NugqSYD6uhGDiRZWqtSJA8g7ihTFNJvVi6kuv4LLt1whHbHCvS8oe7pzP30sfoOjaav9yEi94
NOpa98bUfoZbt/N8x2SLBbqv3ipT2wmG9NkH5Y+vdNXLcLk96fyeRt8Qx8GOL6jBml5timH4ZxdS
QZePAeoLdaDRqSb0CugCCH79iTsOEaNN2BW2PZCceibFBzNlIt1zlNhlcVbnrXlQOA4BysXhy9wg
Tkzm14OBzUx8VFHK6eE6vI1n/20QSEVltAg6HSYqB5YsvSSqgd7ILeCzca2XQqTs0+i3SQHZHsbm
uSHWi9e0TZIhdO3F03DMZrsPYOO9iFlBd1GmOemY+6SBNFKB7/NMTZGdPX+Il/sSrVNlIVtNzbKA
8bT1ZjZBAq01y19oGu1drf0I4bqkvnFwdqy5cnqFgBJiMKhyqTjPRiM+tluEERRKqrnDtJURs9zE
EdK3hwdOPvRjiK8iDpeX2ycd48lbZsBQtDwKUX07+DDnj559+YKnp5hyYO9QY2WwK6ij8mu5sDvx
XRHBxy3R/aFWbYNl3ze4Qtin48ZjyESBitB/h68I/nxlVhHwDsXTf+kzBe/3vqquLOzHu4854zJj
YT/lRuVkIUOAanut/Bi2Xjrodcj27y7xQFfjKVPXuTeshKFfo+ludLZWLYnpxnTXwTF+TxrvGPqy
yBfIf68bCsFX+nHiUuHNjcn2ncrqqOpvv5Zqx3NzNvEDmn30sG6MDUSihHIKwLba8SGk2U5bSNGA
hEVjJNHq6mPl1dhJerHK31ioqJCKTXWgz5zbZUtiiclvrriK24eK9xZJJxog6OQs7qPG5XVnOGMQ
JP3rzfMzU8l/a4pS9l30XKpVEhSIBVy7/s5WuC3Ba8xf1naHjuZXV4gbyqK++PFSAXsxfbyK2tm3
Usas+z7pP9XnUgRubp6yQgUJwfZbUIemER97LRhIh4H62gX/qMQ8hyu8De4HfzepSeGez8+Df9QT
dBx8/SWQqkF+Yjw0ydX9YhN3uLPmQqDLNr4gtAob0duhhs85tnL+/WH50ACuQgPRlpVfAXl0fl2f
Kf8EnKOvnAPxC96C4fLGhanA1EMTXF/qeJz9CeqLiWCXGo1cFL2evHa3/cgkP3+bGXSdFcjGthy2
Yem0DsWN/Fv+7QPomdlc58iYGkMEnDYjBjBFKeRmnuB1m09ngh2kCUsZ2+tm/3KEZGdme2wMAj4p
YqLwCB9nom9Kuc/NlUSBPnfXogbvTxBn8FE76iRDJL0dzZmflhZ8e7kOCMBmQOJMohftTJ4S59J+
vEYn5KRyjhXXOdHGGqMxspA1/Yao4DQh65ZLTtmP9rZ7unCIU0YHimt9spvKgjMq5fdCZtCuz991
DRxA41WvGu9CFoZLxtNcTh3YlwI2MSA9ttsJhw8h1kTFCqmOLo0loTCq3/hEfkgjrYUxG4WQhIHl
WYJPh8J+Ox0by1c7sAIpkKGUinvciAgj/Ryuv1b0hCv3JH/o5cA3zcGkbTpOXZuS2QFy99ZkrAC2
WlHxJCF8aKbs0nPHi6Fhv8tb9lhZK4pzJoXFbSJXTuX7sMr56Q6FNpcXFS0grjMnUjf1lS7QHf3t
mmSlRd+LmuxDBkH6IWlbCrpAhi0w5LbbuLaCRYd9w3fv84bvgXvAJIhaiazYpLhsubgrm7xolMzE
xFw3OmEILDyzyAc3PzrvSEx7w306rxrdEu0CkYr/6b7qwp9MK3BjmJWQGI2nR5ngcEZrbXrpFLSx
kTCHyj7FbeegIWa96WAfw/kOfrVZdGGMeb1PAKFe7yk+NaUk6UAxqIyCDI9i8SOOklPZFJFQvLtn
+8Fa5kULGyCnnadJh13eK0DeuLNXGeuo9yxv75T1zsz06YEasGCaZwsxEb/5C4c6Armpk+66LxqK
3d9irXFb7iHj78Yo9TFv4wR3EJFC9zxYPHODvs7qopuOHNAikgUnSc4huTkXXOvaucVb4bThVPrE
ZMt2WUShyAMlKtC362N6LY0LxyeF4uICuC9VkNjtjeeoIN1ryQG1Vm4QVoibC6dL+Mau/Nx3DDhH
kGJPabL7HT8RLMpjpTc8nmAn0gMolrPbrUHMpbyV5qdrePI0+vuO0dlIxgXY4WvYZNuqGAACVggH
Dbou6HbUHkQRo/xo5wCpUQu7dOMIKc5KAQvXzdH9xF44zc26AQgc3J6/KcpVpIOIUMecPPUNwPk8
BGQRGmGMw0l1A77xsCcoxnGKQn1f8NtNbeFA2bN7/rYAfDzQShwUCZgeaXCkRS6xoxeK17NPnSQW
PffauQQfnpHLGydENpXEVxT6cZgUBFzoAxwVfOeTF4yDgG3BqSvUXcY5Z0zj8DvAWh2iJ1RePU8l
5eZqaI45S6WX1WVcC4A4w2DtkhOICCABz/hvQgAKkvtJ1v8gDaL6G5Y9BqYmlmM6zRNMF+ZDOagJ
qQv9CGQYbmLk9LDnlpiHJRfdp3r7iZpeBEeQBrO78ZQCcY3hIjRGfFuVrINMAWIq2Ta7e0ShJvpR
WIAJ5b2ctHfDeggl7kWXj58c4AryLnwY8QVt7zdfzWSjnztTPrBOXZndOebpA6ibNPuFeKA5zwf6
ooPiYCp2A6O4IPqcgW0JEHv7UV8VxYvVDsZjld6mkaP21If0sVpwZdntL6IuhDszEQ3CPQGYwSov
uAh9CgPVK2Kh0XI73spVPyTSR+WxGcIfxv5sbXTnp5u6TsD9XPOGHqVVSWHD6PcRuG4+bfcT0BYf
LqLNh5Lg2lctOuysTM5Dq3ZQuDOuMh4X8PjLCUP1kV4B4+1GalH8j5DwCBDXTsPzPIvgriDuH9sM
PC9e3TCtmsVEyH7XTXhwqu+dcNzxSgSYP5+OtqWJnf+XNxasncXrPZYfWvoFFzUJTdgbN8Fnd6YD
nQ3lSwhNSJ7U77PNLMJ5uQhOENKSxHcWPYtHnsHnv7EQ2I4EqbNMM+qFGDaDItaaJug30CcpVS2r
PEKI5fcYXhVkr7yHmwAbWVNUgnztlANBTVsf9PLGvLY2Tz9YPZ0+h44Y2Nhf0Tz2R23k8klm7b8S
nIwPHEJkJLG96GvEvJWmliglLGbu25vKtHWruADounOVZQ0fKfdqP7dXJ6YqgMp+ipp1fQlonVZA
d9XTpt0n2HV/3udOBXwpoVWJ8wGtat0JI9qzZ1m/ajUmJFRwLmIBLCzl/KNuBBFu2L3Gyn593koK
tkrTSzldszmw5/DX7pUIHrX6XlRovNYzeC1cXbSCW8EY4prLFmbnR9Z9+5tjJ2Iq6Rp6B+7M4OF3
rdmu+p3u5YnsSU+mi1+nSvPLq9sLAGAmVqleDMpYt/ACNIZZOVTcXQ11wSIBz6vBJaAq3Y3uXboC
68fUMOvvQYq/dT9fQBxZOrLIsZEYStBA8B5p7sQQB4JYw4yy9hPEqhB8cW5utzo4CG9VGCfv6unm
T8GRLUzbHT40gyPuAurvddx6Zbklf2eXy9yQyT5tdShIMFz5tZ5oIi7+siqj0jiJaoOuhuNf7muj
fDVAwuRlcECiJjcc59zeOwmOqDn2CpeayimYrAp2GVTFzhEmTmreWHUs/Mked7G6HyrlgFKRrey2
cKlIeuAGHh6RcEA0eb0JAWw1kQMUPQVFKM8R330eL9vaU6WO3rsCqKxXpbablfCpN/6KQDLXIW8T
zdaUdiHq
`pragma protect end_protected

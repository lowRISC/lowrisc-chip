/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootram (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic         we_i,
   input  logic [63:0]  addr_i,
   input  logic [7:0]   be_i,
   input  logic [63:0]  wdata_i,
   output logic [63:0]  rdata_o
);

   localparam BRAM_SIZE          = 16;        // 2^16 -> 64 KB
   localparam BRAM_WIDTH         = 128;       // always 128-bit wide
   localparam BRAM_LINE          = 2 ** BRAM_SIZE / (BRAM_WIDTH/8);
   localparam BRAM_OFFSET_BITS   = $clog2(64/8);
   localparam BRAM_ADDR_LSB_BITS = $clog2(BRAM_WIDTH / 64);
   localparam BRAM_ADDR_BLK_BITS = BRAM_SIZE - BRAM_ADDR_LSB_BITS - BRAM_OFFSET_BITS;

   initial assert (BRAM_OFFSET_BITS < 7) else $fatal(1, "Do not support BRAM AXI width > 64-bit!");

   // BRAM controller
   wire [7:0] ram_we = we_i ? be_i : 8'b0;

   reg   [BRAM_WIDTH-1:0]         ram [0 : BRAM_LINE-1] = {
128'hf1402973000004933049107300800913, /*    0 */
128'hfe0e9ee3fffe8e9300a00e9311249a63, /*    1 */
128'h00008297011111133ff1011b00004137, /*    2 */
128'h0b42829300008297000280e708e28293, /*    3 */
128'h00000597000280e71305051300000517, /*    4 */
128'h000046b7c10606130000c617fb458593, /*    5 */
128'h240e8e9b000f4eb7011696933ff6869b, /*    6 */
128'hfe0e9ae30085b703fffe8e930005b703, /*    7 */
128'h0006b703ff81011301b111130110011b, /*    8 */
128'h00e6b4230085b70300e6b0230005b703, /*    9 */
128'h00e6bc230185b70300e6b8230105b703, /*   10 */
128'h00000797fcc5cce30206869302058593, /*   11 */
128'h0007806740b787b300d787b301478793, /*   12 */
128'h0000c597305790730907879300000797, /*   13 */
128'h0005b0233bc606130000c617c2458593, /*   14 */
128'h020585930005bc230005b8230005b423, /*   15 */
128'h00100913020004b7017090effec5c6e3, /*   16 */
128'h4009091b02000937004484930124a023, /*   17 */
128'h008979133440297310500073ff24c6e3, /*   18 */
128'h00291913f1402973020004b7fe090ae3, /*   19 */
128'hfe091ee30004a9030009202300990933, /*   20 */
128'hff24c6e34009091b0200093700448493, /*   21 */
128'hffdff06f1050007334102373342022f3, /*   22 */
128'h6e61697241206d6f7266206f6c6c6548, /*   23 */
128'h61207469617720657361656c50202165, /*   24 */
128'h00000000000a2e2e2e746e656d6f6d20, /*   25 */
128'h00000000000000000000000000000000, /*   26 */
128'h00000000000000000000000000000000, /*   27 */
128'h00000000000000000000000000000000, /*   28 */
128'h00000000000000000000000000000000, /*   29 */
128'h00000000000000000000000000000000, /*   30 */
128'h00000000000000000000000000000000, /*   31 */
128'hd963454c0005cc635735c28587ae6914, /*   32 */
128'he21c97b6470102a787b30a00051300b7, /*   33 */
128'h853e85b200030563018533038082853a, /*   34 */
128'h8f8686930000c697b7edfda007138302, /*   35 */
128'h87930000c7976294a24707130000c717, /*   36 */
128'h87b30280069302d787bb878d8f99a1a7, /*   37 */
128'h47148082853a470100e7956397ba02d7, /*   38 */
128'hf0efe4061141b7f502870713fea68de3, /*   39 */
128'hbfe545018082014160a26108c509fbbf, /*   40 */
128'hf0efe852ec4ef04af426f822fc067139, /*   41 */
128'h0000ba17440144814985892acd31f9bf, /*   42 */
128'hc091553500f44d6300c9278347ca0a13, /*   43 */
128'h61216a4269e2790274a2744270e24501, /*   44 */
128'h67a2ed19f29ff0ef854a85a200308082, /*   45 */
128'h50ef8552000995632485cb990087c783, /*   46 */
128'h0513bf652405230080ef498165224ae0, /*   47 */
128'hf2dff0efe42ef406f0227179b7c1fda0, /*   48 */
128'h842aee7ff0ef083065a2c105fda00413, /*   49 */
128'h00f7096300c547030ff007936562e911, /*   50 */
128'h547980826145740270a285221f6080ef, /*   51 */
128'hf0efec4ef04af426f822fc067139bfd5, /*   52 */
128'h0000a9970ff00913440184aacd01eebf, /*   53 */
128'h74a2744270e200f4496344dc59498993, /*   54 */
128'hf0ef852685a200308082612169e27902, /*   55 */
128'h85a20127896300c7c78367a2ed09e83f, /*   56 */
128'hb7d92405190080ef652240a050ef854e, /*   57 */
128'he8dff0ef892eec26f406e84af0227179, /*   58 */
128'he45ff0ef84aa85ca0030c11dfda00413, /*   59 */
128'h538505130000a517864a608ced01842a, /*   60 */
128'h740270a28522152080ef65223cc050ef, /*   61 */
128'hf406ec26f022717980826145694264e2, /*   62 */
128'h85a6842ac11dfda00413e47ff0ef84ae, /*   63 */
128'hcf63445c394050ef510505130000a517, /*   64 */
128'h5435118080ef50e505130000a51700f4, /*   65 */
128'h003085228082614564e2740270a28522, /*   66 */
128'h0ec080ef6522f565842adcfff0ef85a6, /*   67 */
128'h5479fcf71be30ff0079300c7c70367a2, /*   68 */
128'he50965a2de1ff0eff406e42e7179bfc1, /*   69 */
128'hf96dd97ff0ef08308082614570a24501, /*   70 */
128'he42eec064108842ae8221101bfc56562, /*   71 */
128'h852200030e6302053303c919db9ff0ef, /*   72 */
128'h60e2fda005138302610560e265a26442, /*   73 */
128'h0000b7977139bfdd4501808261056442, /*   74 */
128'h04130000b417f426f822639c68478793, /*   75 */
128'h043b840d8c057a2484930000b4977aa4, /*   76 */
128'h892afc06e852ec4ef04a0280079302f4, /*   77 */
128'h942602f4043344ea0a130000aa1789ae, /*   78 */
128'h69e2790274a2744270e2450100849b63, /*   79 */
128'h290050ef855285ca6090808261216a42, /*   80 */
128'hbfc902848493c50169d060ef854a608c, /*   81 */
128'hb7e16522f569cdbff0ef852685ce0030, /*   82 */
128'h84b68432e42efc06f04af426f8227139, /*   83 */
128'hcb5ff0ef083065a2c115cf7ff0ef893a, /*   84 */
128'h70e2978285a2615c862686ca6562e519, /*   85 */
128'hbfc5fda0051380826121790274a27442, /*   86 */
128'h84b68432e42efc06f04af426f8227139, /*   87 */
128'hc75ff0ef083065a2c115cb7ff0ef893a, /*   88 */
128'h70e2978285a2655c862686ca6562e519, /*   89 */
128'hbfc5fda0051380826121790274a27442, /*   90 */
128'hc7dff0ef84b2e42ef822fc06f4267139, /*   91 */
128'h701ce509c39ff0ef842a083065a2c105, /*   92 */
128'h8082612174a2744270e2978285a66562, /*   93 */
128'h2785c3190017f713419cbfcdfda00513, /*   94 */
128'hd71b8e5927a106220086571b419cc19c, /*   95 */
128'h0ff77713c19c0087d7138ed906a20086, /*   96 */
128'h122300d5112300c510238fd90087979b, /*   97 */
128'hf022f4067179419c80820005132300f5, /*   98 */
128'h419c00f510230457879b6785c19c27d1, /*   99 */
128'h0087979b0ff777130087d713c632842a, /*  100 */
128'hc4360509084c57fd460900f11a238fd9, /*  101 */
128'h051301610593460978b060ef00f11b23, /*  102 */
128'h00041323082c462147c177d060ef0044, /*  103 */
128'h00f404a347c5769060efec3e00840513, /*  104 */
128'h753060ef00c4051300041523006c4611, /*  105 */
128'h01440693747060ef01040513002c4611, /*  106 */
128'hfed79ce39f31ffe7d6030789470187a2, /*  107 */
128'h9fb94107d71b9fb9934117424107579b, /*  108 */
128'h80826145740270a200f41523fff7c793, /*  109 */
128'h97ba46a167856398538787930000b797, /*  110 */
128'hc7bb27850077e793fff6079b8007bc23, /*  111 */
128'h3823973e678500f547636805450102d7, /*  112 */
128'h010686bb0035169b0005b883808280c7, /*  113 */
128'he0221141bff105a125050116b02396ba, /*  114 */
128'hfa5ff0efe406450185aa86220005841b, /*  115 */
128'hec26f022717980820141640260a28522, /*  116 */
128'h693060efe436f4064619051984b2842a, /*  117 */
128'h162347a1687060ef85b64619852266a2, /*  118 */
128'h614564e200e4859b70a27402852200f4, /*  119 */
128'h3a8130236785737dc5010113fadff06f, /*  120 */
128'h3931342338913c233a11342339213823, /*  121 */
128'h377134233761382337513c2339413023, /*  122 */
128'h3507879335a1382335913c2337813023, /*  123 */
128'hce042023d00007b7943e747d978a911a, /*  124 */
128'hd0040023f0040023e0040023ca040b23, /*  125 */
128'ha51785aa00e7ea63892a5800073797aa, /*  126 */
128'h00054703a0017a7040ef152505130000, /*  127 */
128'h970a3507871374fd678526f711634789, /*  128 */
128'hcb848b13970a350787139abacd848a93, /*  129 */
128'h9c3a9b3a49818a368cb28baed0048c13, /*  130 */
128'hc7830015cd03013907b395ca0f098593, /*  131 */
128'h869b01a989bb058902a0071329890f07, /*  132 */
128'h24e78163471904f76b6326e78d630007, /*  133 */
128'hcc848513470d2ae78963470502f76263, /*  134 */
128'h40ef252505130000a51785b622e78963, /*  135 */
128'hfee794e3473d22e785634731b77d71f0, /*  136 */
128'h953e866ae0048513978a350787936785, /*  137 */
128'h03600713b759e00d002354d060ef9d22, /*  138 */
128'h22e780630330071300f76e6322e78363, /*  139 */
128'haad94605cb648513fae798e303500713, /*  140 */
128'hf8e79ce30ff0071324e7856303800713, /*  141 */
128'h24e781630007859b747d471500614783, /*  142 */
128'h000ca7833ae79d63470938e781634719, /*  143 */
128'h05134985978a350a87936a8516079263, /*  144 */
128'h60ef013ca023953e461101090593ce44, /*  145 */
128'h01490593ce840513978a350a87934d10, /*  146 */
128'h028505130000a5174bb060ef953e4611, /*  147 */
128'h978a350a8793657040efde0254e25a52, /*  148 */
128'h441060ef854a55fd4619993ecf840913, /*  149 */
128'h879346f115231350079300f103a3478d, /*  150 */
128'h85a6460594becb740493c2a6978a350a, /*  151 */
128'h06a303200793469060efc0d246c10513, /*  152 */
128'h4a1195becf040593978a350a879346f1, /*  153 */
128'h0793445060ef4741072346f105134611, /*  154 */
128'hcf440593978a350a879346f109a30360, /*  155 */
128'h423060ef47410a2347510513461195be, /*  156 */
128'h03a346f10ca347b1051385a6460557fd, /*  157 */
128'h061310200793409060ef47310d230001, /*  158 */
128'h07933a3060efde3e37a1051345810f00, /*  159 */
128'h3961051385de4799464136f11d231010, /*  160 */
128'h13232637879377e13db060ef36f10e23, /*  161 */
128'h350a879346f1142335378793679946f1, /*  162 */
128'h0440061304300693943ecec40413978a, /*  163 */
128'h85a2460156fdba1ff0ef3721051385a2, /*  164 */
128'h0e8885de86ca5672bd5ff0ef35e10513, /*  165 */
128'h3a0134033a813083911a6305cebff0ef, /*  166 */
128'h38013a03388139833901390339813483, /*  167 */
128'h36013c0336813b8337013b0337813a83, /*  168 */
128'h851380823b01011335013d0335813c83, /*  169 */
128'ha00d953e978a3507879367854611cd04, /*  170 */
128'h953e866af0048513978a350787936785, /*  171 */
128'h85564611b39df00d002332d060ef9d22, /*  172 */
128'h87936785bfdd855a4611bbb131f060ef, /*  173 */
128'h303060ef4611953ece048513978a3507, /*  174 */
128'h00f40123ce14478300f401a3ce044783, /*  175 */
128'h00f40023ce34478300f400a3ce244783, /*  176 */
128'h866ab759cc048513bb29cef42023401c, /*  177 */
128'h2783b311d00d00232cb060ef9d228562, /*  178 */
128'h0000a51700fa2023478512079a63000a, /*  179 */
128'h0e88010905934611459040efe3c50513, /*  180 */
128'hcb840513978a35048793648529f060ef, /*  181 */
128'h35314703287060ef014905934611953e, /*  182 */
128'h0000a517350145833511460335214683, /*  183 */
128'h00a1468335015783419040efe0c50513, /*  184 */
128'h352157831cf71e230000b71700914603, /*  185 */
128'h0000b717e0c505130000a51700814583, /*  186 */
128'h01b147033e5040ef00b147031cf71323, /*  187 */
128'h0000a517018145830191460301a14683, /*  188 */
128'h01214683013147033c9040efe0c50513, /*  189 */
128'he10505130000a5170101458301114603, /*  190 */
128'h05130000a51755c2010157833ad040ef, /*  191 */
128'hb7170121578316f713230000b717e1e5, /*  192 */
128'hf6bb02f5d63b03c0079314f71e230000, /*  193 */
128'h02f5d5bbe107879b678502f6763b02f5, /*  194 */
128'h95bee0040593978a3504879336d040ef, /*  195 */
128'h35048793355040efdf8505130000a517, /*  196 */
128'hdf0505130000a51795be978af0040593, /*  197 */
128'h40efdfa505130000a517b50133d040ef, /*  198 */
128'h20234785de0796e3000a2783bbcd32f0, /*  199 */
128'ha517313040efdee505130000a51700fa, /*  200 */
128'h350787936785307040efdf2505130000, /*  201 */
128'hdf8505130000a51795be978ad0040593, /*  202 */
128'hb35d2e3040efdfe505130000a517bf45, /*  203 */
128'hf852fc4ee0cae4a6e8a2ec86711d737d, /*  204 */
128'h6a85e12505130000a517911a89aaf456, /*  205 */
128'h0493978a020a8793747d2bb040efca02, /*  206 */
128'hb7970a3060ef852655fd461994beff84, /*  207 */
128'hc83e4a05fef40913439cf02787930000, /*  208 */
128'h993e978a020a879312f11d2313500793, /*  209 */
128'h07930c5060ef014107a31a68460585ca, /*  210 */
128'h020a879312f10f23479112f10ea30370, /*  211 */
128'h60ef13f10513461195beff040593978a, /*  212 */
128'h14f101a314510513460585ca57fd0a10, /*  213 */
128'h0fc00793087060ef000107a315410223, /*  214 */
128'h021060efca3e04a1051345810f000613, /*  215 */
128'h05134641479985ce04f1152310100793, /*  216 */
128'h2637879377e1059060ef04f106230661, /*  217 */
128'h879312f11c2335378793679912f11b23, /*  218 */
128'h06930421051385a2943e1451978a020a, /*  219 */
128'h02e1051385a2821ff0ef044006130430, /*  220 */
128'h85ce86a610084652855ff0ef460156fd, /*  221 */
128'h64a66446450160e6911a630596bff0ef, /*  222 */
128'ha51785aa808261257aa27a4279e26906, /*  223 */
128'h3423810101131970406fd02505130000, /*  224 */
128'h34237d2138237c913c237e8130237e11, /*  225 */
128'h893689b2e04605a1051384aa71597d31, /*  226 */
128'h101867857b6060efd602e83eec3ae442, /*  227 */
128'h943e7fc404136762747d97ba81078793, /*  228 */
128'hf8aff0efd64e0521051385a2864a86ba, /*  229 */
128'hf0ef03e10513863e86c285a267c26822, /*  230 */
128'h8cfff0ef86c685a6180856326882fbaf, /*  231 */
128'h7d8134837e01340345017e8130836165, /*  232 */
128'h716d80827f0101137c8139837d013903, /*  233 */
128'h003547830045480300554883e222e606, /*  234 */
128'ha597842a000546030015468300254703, /*  235 */
128'h40efc52505130000a517c52585930000, /*  236 */
128'ha597860ac10d842adedff0ef85220cf0, /*  237 */
128'h40efc5a505130000a517c32585930000, /*  238 */
128'h0000a51780826151641260b285220af0, /*  239 */
128'h091040efde07ae230000b797c7450513, /*  240 */
128'hf85afc56e0d2e4ceeca6f0a27159b7cd, /*  241 */
128'h8a2ae46ee8caf486e86aec66f062f45e, /*  242 */
128'h918a8a930000ba974401ff05049389ae, /*  243 */
128'h0000ac1706000b93c48b0b130000ab17, /*  244 */
128'hfff58d1bc44c8c930000ac97c54c0c13, /*  245 */
128'h6a0669a6694664e6740670a603344163, /*  246 */
128'h61656da26d426ce27c027ba27b427ae2, /*  247 */
128'h011040ef855ae7a9c42900f477938082, /*  248 */
128'hfe05879b0007c583012487b34dc14901, /*  249 */
128'h09057f2040ef856602fbe2630ff7f793, /*  250 */
128'h7e0040ef774505130000a517ffb912e3, /*  251 */
128'hb7c57d2040ef8562a0317da040ef8556, /*  252 */
128'h40efbd2505130000a5170104c583dbe5, /*  253 */
128'h00f979134d81fffd4913028d1d637be0, /*  254 */
128'h855aff2dcce32d857a8040ef8556a029, /*  255 */
128'h00f45b630009079bff04791379c040ef, /*  256 */
128'h04852405784040ef718505130000a517, /*  257 */
128'hf793fe05879b0007c583012a07b3b781, /*  258 */
128'hb7e90905764040ef856600fbe7630ff7, /*  259 */
128'he44ee84aec267179bfdd75a040ef8562, /*  260 */
128'h86930000a697893289ae84b6f022f406, /*  261 */
128'h00009717b4c686930000a697c50939e6, /*  262 */
128'h854a85a6b44606130000a617ffc70713, /*  263 */
128'h85bb00955d6300098f63842a6dc040ef, /*  264 */
128'h40ef954ab2c606130000a61786ce40a4, /*  265 */
128'hffd4841b00f44463ffe4879b9c296be0, /*  266 */
128'h276060efafc585930000a59700890533, /*  267 */
128'h8082614569a2694264e2854a740270a2, /*  268 */
128'h0613002c7115f73ff06f4581862e86b2, /*  269 */
128'h0000a517002cfebff0efed8645050c80, /*  270 */
128'h8082612d450160ee6a8040efae450513, /*  271 */
128'h47b704a76963862e9ff787133b9ad7b7, /*  272 */
128'hf7633e70079304a7676323f78713000f, /*  273 */
128'hae8707130000b7173e80079346890ca7, /*  274 */
128'he426e822ec0600074903e04a97361101, /*  275 */
128'ha51785aa690264a260e2644202091663, /*  276 */
128'h879346816440406f6105a8a505130000, /*  277 */
128'h02f57433bf7d240787934685b7d9a007, /*  278 */
128'h0287e66347293e800793c02102f555b3, /*  279 */
128'h0287746306300713c70502f4773347a9, /*  280 */
128'h0324341302e4743302f457b306400713, /*  281 */
128'h5433bfc102e45433a039943e00144413, /*  282 */
128'h40ef84b2a34505130000a517f86102f4, /*  283 */
128'h40efa2a505130000a51785a2c8015de0, /*  284 */
128'ha517690264a285ca862660e264425ce0, /*  285 */
128'ha51785aa5b40406f6105a1a505130000, /*  286 */
128'h481958d94781862eb78d9ea505130000, /*  287 */
128'h1782cd8500e555b303c6871b02f886bb, /*  288 */
128'he42697c211019f6808130000b8179381, /*  289 */
128'h60e26442e495e04ae822ec060007c483, /*  290 */
128'h61059ca505130000a51785aa690264a2, /*  291 */
128'h0000a51785aafb079de3278555c0406f, /*  292 */
128'hfff7c79300e797b357fdb7f59b450513, /*  293 */
128'h03b6869b02f5053347a9c10d44018d7d, /*  294 */
128'hf46300e45433942a47a500d414334405, /*  295 */
128'h8932962505130000a517058514590087, /*  296 */
128'h958505130000a51785a2c80150c040ef, /*  297 */
128'h64a2690285a6864a60e264424fc040ef, /*  298 */
128'h71514e20406f6105960505130000a517, /*  299 */
128'he96ae5cee9caf1a202c7073b8cbaed66, /*  300 */
128'he56ef162f55ef95afd56e1d2eda6f586, /*  301 */
128'h00e7f66384368d3289ae892a04000793, /*  302 */
128'hdcbb4cc1000c956302ccdcbb04000c93, /*  303 */
128'h0017849be03e020d1a13001d179b03ac, /*  304 */
128'h908b0b130000ab1703810a93020a5a13, /*  305 */
128'h7d8c0c1300008c17870b8b930000ab97, /*  306 */
128'h6a0e69ae694e64ee740e70ae4501e00d, /*  307 */
128'h616d6daa6d4a6cea7c0a7baa7b4a7aea, /*  308 */
128'h440040ef8c4505130000a51785ca8082, /*  309 */
128'h470186ce000c8d9b008cf46300040d9b, /*  310 */
128'h971305b66c630007061b430948a14811, /*  311 */
128'h06bb0d9de66399ba034707339301020d, /*  312 */
128'h415705bb0006861b02e00813875603bd, /*  313 */
128'h05130000a51785d6963e011c0ac5ed63, /*  314 */
128'h043b66a23e4040effa060c23e43687e5, /*  315 */
128'h557dd1350c0070ef99369281168241b4, /*  316 */
128'h260195d6002715934290030d1b63b795, /*  317 */
128'hec42f046f41a855a658292011602c190, /*  318 */
128'h96d27322674266a23a8040efe436e83a, /*  319 */
128'h15936290011d1863bf85686278820705, /*  320 */
128'h0006d603006d1c63bfc1e19095d60037, /*  321 */
128'hbf6500c590239241164295d600171593, /*  322 */
128'h00c580230ff6761300ea85b30006c603, /*  323 */
128'h6ae3270567220ec070efe43a855eb75d, /*  324 */
128'h053300074583bfdd4701bf1d3cfdfe97, /*  325 */
128'h0185959bc519097575130005450300bc, /*  326 */
128'hbf390705010700230005d4634185d59b, /*  327 */
128'h8082e21c00b7f4634501918187aa1582, /*  328 */
128'h89aa04000613fd4e7115bfd58f8d2505, /*  329 */
128'hf556f952e1cae5a6e9a2ed8600884581, /*  330 */
128'h577d67869982e16ae566e962ed5ef15a, /*  331 */
128'h55796318674707130000a7178ff98361, /*  332 */
128'h00009b174a8503800a13440106e79d63, /*  333 */
128'h80000c3778cb8b9300009b97754b0b13, /*  334 */
128'h07815783764d0d1300009d1708000cb7, /*  335 */
128'h06137786028a05bba091656600f46463, /*  336 */
128'h77c20957926347a299829dbd00280380, /*  337 */
128'h040908637922276040ef855a85a2cfbd, /*  338 */
128'h0000951785a60397e863018487b37482, /*  339 */
128'h64ae644e60ee5575258040ef70450513, /*  340 */
128'h6caa6c4a6bea7b0a7aaa7a4a79ea690e, /*  341 */
128'h40ef856a86ca85a666428082612d6d0a, /*  342 */
128'h77a274c2998285260009061b45c222e0, /*  343 */
128'h855e85ca993e86268c9d79020097ff63, /*  344 */
128'h2405002060ef854a4581862620c040ef, /*  345 */
128'ha7178082400005378082057e4505bfb1, /*  346 */
128'h869300756513157d631c77a707130000, /*  347 */
128'h057e450597aa20000537e30895360017, /*  348 */
128'h862a0ce507638207871367858082953e, /*  349 */
128'h6b050513000095178087871308a74463, /*  350 */
128'h000095178006079b04c7496306e60b63, /*  351 */
128'h0000951787f787936785c3ad68c50513, /*  352 */
128'h11417c07879b77fd04c7c96370c50513, /*  353 */
128'h05130000a5176fe58593000095979e3d, /*  354 */
128'h05130000a51760a2144040efe4066de5, /*  355 */
128'h05130000951781078713808201416ce5, /*  356 */
128'h0513000095178187879300e60a6365e5, /*  357 */
128'h00009517830787138082faf612e365e5, /*  358 */
128'h8287879300c74963fee609e367c50513, /*  359 */
128'h951783878713bfe96585051300009517, /*  360 */
128'h951784078793fce608e366a505130000, /*  361 */
128'h6205051300009517bf7566a505130000, /*  362 */
128'h84ae892af406e84aec26f02271798082, /*  363 */
128'h942a9041144201045513029044634401, /*  364 */
128'h1542fff54513740270a2952201045513, /*  365 */
128'h0068460985ca808261459141694264e2, /*  366 */
128'h00f107a334f9090900c147836ff050ef, /*  367 */
128'hbf55943e00e1578300f1072300d14783, /*  368 */
128'h8793f44ef84afc26e486e0a26785715d, /*  369 */
128'h0e636dd7879367a13cf50563842e8067, /*  370 */
128'h082884b205e944079a638005079b0af5, /*  371 */
128'ha517461985ca006409136ad050ef4611, /*  372 */
128'h079301744583699050ef5d2505130000, /*  373 */
128'h1cf5826347b108b7e76332f5896302e0, /*  374 */
128'h478502b7e3631af58363479104b7e563, /*  375 */
128'h83635aa5051300009517478910f58463, /*  376 */
128'ha41d002040ef746505130000951702f5, /*  377 */
128'h5b0505130000951747a118f582634799, /*  378 */
128'h2cf5826347f5a4317e9030effef591e3, /*  379 */
128'h0000951747d916f58a6347c500b7ed63, /*  380 */
128'h866302100793bf6dfef580e35cc50513, /*  381 */
128'h051300009517faf596e3029007932af5, /*  382 */
128'h04b7e2632cf5826306200793b7c95e65, /*  383 */
128'h02f0079300b7ef632af5826303300793, /*  384 */
128'h5e850513000095170320079328f58763, /*  385 */
128'h079328f5846305c00793b7bdf8f58ae3, /*  386 */
128'hbf91f6f58de35fe505130000951705e0, /*  387 */
128'h0670079300b7ef6328f5866308400793, /*  388 */
128'h610505130000951706c0079326f58b63, /*  389 */
128'h079326f5886308900793b73df4f58ae3, /*  390 */
128'h9517f0f59ce30880079326f589630ff0, /*  391 */
128'h0000a79701e45703b73d61a505130000, /*  392 */
128'h12f714634dc989930000a9974e47d783, /*  393 */
128'h10f71c634ce7d7830000a79702045703, /*  394 */
128'h0000a5974619539050ef852285ca4619, /*  395 */
128'h012301a45783529050ef854a49c58593, /*  396 */
128'h859b01c4578300f41f23020412230204, /*  397 */
128'h1d230009d78302f4102302240513fde4, /*  398 */
128'h0ea3db9ff0ef00f41e230029d78300f4, /*  399 */
128'h1223862601c1578300a10e23812100a1, /*  400 */
128'h00009517a06ddcbfe0ef450185a202f4, /*  401 */
128'hb55942a5051300009517bd4141c50513, /*  402 */
128'h470302444783bdb54385051300009517, /*  403 */
128'h178300f10e230254478300f10ea30264, /*  404 */
128'h00e10e2327810274470300e10ea301c1, /*  405 */
128'h0234470300e10ea301c1190302244703, /*  406 */
128'h04e79b6301c156830450071300e10e23, /*  407 */
128'h0000a597461947e23ad79e230000a797, /*  408 */
128'h0000a71739c505130000a51739458593, /*  409 */
128'ha79766a24762449050efe43638f72e23, /*  410 */
128'h450102a40593ff89061b372787930000, /*  411 */
128'h616179a2794274e2640660a655a060ef, /*  412 */
128'h0000a71747e204e69463043007138082, /*  413 */
128'hc799439c360787930000a79734f72e23, /*  414 */
128'h0000a697f7e9439c350787930000a797, /*  415 */
128'h0000a597340606130000a61734468693, /*  416 */
128'h0713b765d6dfe0ef02a4051334458593, /*  417 */
128'h30ef352505130000951702e798634d20, /*  418 */
128'h051300009517cdcff0ef852285a656f0, /*  419 */
128'hcc6ff0ef02a4051385ca55b030ef34e5, /*  420 */
128'h67c101e45703f6e787e35fe00713bf95, /*  421 */
128'h4611f4f70de302045703f6f701e317fd, /*  422 */
128'hb799375050ef0868300585930000a597, /*  423 */
128'h051300009517b3353285051300009517, /*  424 */
128'h9517bb213445051300009517b30d32e5, /*  425 */
128'h3685051300009517b339352505130000, /*  426 */
128'h00009517b9ed36e5051300009517b311, /*  427 */
128'hb1dd39a5051300009517b9c538c50513, /*  428 */
128'h051300009517b9f13b05051300009517, /*  429 */
128'hd703b1e13e45051300009517b9c93d65, /*  430 */
128'h84930000a49727e7d7830000a7970265, /*  431 */
128'hd7830000a7970285d703ecf711e32764, /*  432 */
128'h89930205891320000793eaf719e32687, /*  433 */
128'h2c3050ef854a85ce461900f59a230165, /*  434 */
128'h2b3050ef854e226585930000a5974619, /*  435 */
128'h50ef00640513216585930000a5974619, /*  436 */
128'h01c45783297050ef852285ca46192a10, /*  437 */
128'h02f4142301e4578302f4132302a00613, /*  438 */
128'h00f41f230024d78300f41e230004d783, /*  439 */
128'h0000951785aab36900f4162360800793, /*  440 */
128'h430017b7bba54601409030ef36c50513, /*  441 */
128'h74132601608130239f0101138307b603, /*  442 */
128'h8406871b0387759366850034171b00f6, /*  443 */
128'h3c23630c8387b783972a430005379f2d, /*  444 */
128'h5f200813ffc5849b2581601134235e91, /*  445 */
128'h00c5963b101005938a1d08b8696335b9, /*  446 */
128'h87930000a797cfb527818ff1fff7c793, /*  447 */
128'h869b7007f7930084179bea25439014e7, /*  448 */
128'h00d100a3872646d496aa068e9ebd8006, /*  449 */
128'h00d100230086d69b0106d69b0106969b, /*  450 */
128'h806686936685c6918005069b00015503, /*  451 */
128'h67139fad377d8005859b658502d51a63, /*  452 */
128'h868a83f502d7473b1782270546a10077, /*  453 */
128'h862602e6446397c285b6430008378f95, /*  454 */
128'h30838287b823430017b70405aa1ff0ef, /*  455 */
128'h610101135f8134838526600134036081, /*  456 */
128'hbc2306a126050008380300d788338082, /*  457 */
128'he42643c0e8220c2007b71101b7e1ff06, /*  458 */
128'h16938304b703430014b747812401ec06, /*  459 */
128'h2485051300009517e7990206c1630337, /*  460 */
128'h64a2644260e2c3c00c2007b72cd030ef, /*  461 */
128'hf0227179bfc14785eb9ff0ef80826105, /*  462 */
128'h078585930000a597461184ae8432ec26, /*  463 */
128'h030787930000a7970eb050eff4060068, /*  464 */
128'h88930000a89785a6862247b20007a803, /*  465 */
128'ha5170450069301a757030000a7170168, /*  466 */
128'h740270a285228d4ff0ef022505130000, /*  467 */
128'h15428d5d05220085579b8082614564e2, /*  468 */
128'h8fd966c10185579b0185171b80829141, /*  469 */
128'h0085151b8fd98f750085571bf0068693, /*  470 */
128'h07b7715d808225018d5d8d7900ff0737, /*  471 */
128'hc63e04b0051345854601007427f90900, /*  472 */
128'h70efec56f052f44efc26e0a2f84ae486, /*  473 */
128'h1f1030ef1845051300009517892a0770, /*  474 */
128'h57b90a091d63c31901079713fff94793, /*  475 */
128'h03a30000a7175785f8f708230000a717, /*  476 */
128'ha717578df6f70f230000a7175789f8f7, /*  477 */
128'hf6f706230000a7175791f6f70aa30000, /*  478 */
128'h8da30000a797fe056513893d003070ef, /*  479 */
128'h50ef0048f4e585930000a5974611f4a7, /*  480 */
128'h50ef0028f3c585930000a59746097e00, /*  481 */
128'h0613010006374722f31ff0ef45127d00, /*  482 */
128'h15020ff777138ff183210087179bf006, /*  483 */
128'h93c180a6b02317c29101430016b78fd9, /*  484 */
128'h640660a68086b7838006b78380f6b423, /*  485 */
128'h6ae27a0279a2794274e282f6b42347a1, /*  486 */
128'h8a930000aa9744010280049380826161, /*  487 */
128'h0099563349990b6a0a1300009a17ed6a, /*  488 */
128'h00c780230004059b0ff67613015407b3, /*  489 */
128'hbf91ff3411e334e10f9030ef04058552, /*  490 */
128'h073771398087b5838007b603430017b7, /*  491 */
128'hf04af426f822fc068f4d91c115c20080, /*  492 */
128'h0000951780e7b423e05ae456e852ec4e, /*  493 */
128'he6b747030000a7170b9030ef07450513, /*  494 */
128'he5d848030000a817e647c7830000a797, /*  495 */
128'he49646030000a617e526c6830000a697, /*  496 */
128'h0485051300009517e405c5830000a597, /*  497 */
128'h00044783e2c404130000a41707d030ef, /*  498 */
128'h0f230000a717e06989930000a9974481, /*  499 */
128'h6a89dfaa0a130000aa1700144783e0f7, /*  500 */
128'h00262b3700244783e0f704a30000a717, /*  501 */
128'h00344783def70b230000a71743001937, /*  502 */
128'h0000a71700444783def705a30000a717, /*  503 */
128'hdcf70aa30000a71700544783def70023, /*  504 */
128'hda07a0230000a797da0796230000a797, /*  505 */
128'hd807ae230000a797da07a4230000a797, /*  506 */
128'he78d0009a783e4a9d807a8230000a797, /*  507 */
128'h9713830937835a0b0493eddfe0ef8522, /*  508 */
128'h5de30337971383093783020745630337, /*  509 */
128'hdff154fd000a2783bfc5bbbff0effc07, /*  510 */
128'hba1ff0efbfc1710a849377d050ef4501, /*  511 */
128'h07a20005470300154783b7d914fdb7e9, /*  512 */
128'h05628fd907c200354503002547838f5d, /*  513 */
128'h808200f61363367d57fd808225018d5d, /*  514 */
128'h57fdb7f5fee50fa3058505050005c703, /*  515 */
128'hbfcd050500b50023808200f61363367d, /*  516 */
128'h00958413e04ae426ec06e8221101495c, /*  517 */
128'h481586ca02000513478101853903cfa5, /*  518 */
128'h0e6327850006c703462d02e0031348a5, /*  519 */
128'h0023011795630e5007130107146300a7, /*  520 */
128'hfcc79ee30685040500e4002304050064, /*  521 */
128'hf0ef00f5842384ae01c9051300b94783, /*  522 */
128'h0087979b0189470301994783c088f59f, /*  523 */
128'h979b016947030179478300f492238fd9, /*  524 */
128'h644260e20004002300f493238fd90087, /*  525 */
128'h0593cf99873e611c80826105690264a2, /*  526 */
128'h986302d5fc630007468303a006130200, /*  527 */
128'h0705a00d577d00d706630017869300c6, /*  528 */
128'hf593fd06869b577d46050007c683b7dd, /*  529 */
128'h853ae11c0006871b078900b666630ff6, /*  530 */
128'h611cc915bfd5c56747030000a7178082, /*  531 */
128'h008557030067d683c70d0007c703cb85, /*  532 */
128'h3c4060ef0017c503e406114102e69063, /*  533 */
128'h8082014160a24525c391450100157793, /*  534 */
128'h979b468d01a5c70301b5c78380824525, /*  535 */
128'h0155c78300d51d630007079b8f5d0087, /*  536 */
128'h8fd90107979b8fd50087979b0145c683, /*  537 */
128'h5904e44eec26f02271798082853e2781, /*  538 */
128'h00154503842a03450993e052e84af406, /*  539 */
128'h505ce1312501352060ef85ce86264685, /*  540 */
128'h450100e7eb6340f487bb000402234c58, /*  541 */
128'h808261456a0269a2694264e2740270a2, /*  542 */
128'h001445034c5cff2a74e34a0500344903, /*  543 */
128'hb7e5397d310060ef85ce86269cbd4685, /*  544 */
128'h4501f8dff06fc39900454783b7f94505, /*  545 */
128'h4401e04ae426ec06e8221101591c8082, /*  546 */
128'h0005041bfddff0ef892e84aa02b78763, /*  547 */
128'h60ef03448593864a46850014c503ec19, /*  548 */
128'h85220324a823597d4405c11925012980, /*  549 */
128'he822110180826105690264a2644260e2, /*  550 */
128'h842ad91c0005022357fde04ae426ec06, /*  551 */
128'h2324470323344783e52d2501fa3ff0ef, /*  552 */
128'hd79b776d0107979b8fd90087979b4509, /*  553 */
128'hf0ef06a4051302f71f63a55707134107, /*  554 */
128'h4537fff50913010005370005079bd59f, /*  555 */
128'h00978c6345010127f7b3146504930054, /*  556 */
128'h8d05012575332501d33ff0ef08640513, /*  557 */
128'h80826105690264a2644260e200a03533, /*  558 */
128'hfc26e0a2e486f44ef84a715dbfcd450d, /*  559 */
128'h8932852e89aa00053023e85aec56f052, /*  560 */
128'ha7970035171302054e6347addd9ff0ef, /*  561 */
128'hc01547b184aa638097baa5a787930000, /*  562 */
128'h60ef00144503cb85000447830089b023, /*  563 */
128'hc111891100090563e38d001577931e20, /*  564 */
128'h6ae27a0279a2794274e2640660a647a9, /*  565 */
128'h000400230ff4f51380826161853e6b42, /*  566 */
128'hfb71478d001577130f4060ef00a400a3, /*  567 */
128'hee1ff0ef85224581f569891100090463, /*  568 */
128'h23a40a131fa40913848a04f51a634785, /*  569 */
128'hc5bff0ef854ac7894501ffc9478389a6, /*  570 */
128'h8913ff2a14e30991094100a9a0232501, /*  571 */
128'h852285d6000a876345090004aa830104, /*  572 */
128'h4785470dfe9915e30491c10de9dff0ef, /*  573 */
128'h4a81f6e504e34785470db7bd00e51963, /*  574 */
128'h979b03f4470304044783bfb947b5c119, /*  575 */
128'h200007134107d79b0107979b8fd90087, /*  576 */
128'h0089999b04a4478304b44983fef711e3, /*  577 */
128'h2e230444490329811a09866300f9e9b3, /*  578 */
128'h0ff7f793012401a3fff9079b47050134, /*  579 */
128'hfa0b03e30164012304144b03faf769e3, /*  580 */
128'h478304644a03ffc900fb77b3fffb079b, /*  581 */
128'h77930144142300fa6a33008a1a1b0454, /*  582 */
128'h0085151b0474448304844503f3c100fa, /*  583 */
128'h2501042447030434478314050e638d45, /*  584 */
128'h571b2781033906bbdfb18fd90087979b, /*  585 */
128'h04bbf4c564e3873200d7063b9f3d004a, /*  586 */
128'h664119556905dd8d84ae0364d5bb40c5, /*  587 */
128'h873b490d00b673630905165500b93933, /*  588 */
128'h03542023cc04d458015787bb248900ea, /*  589 */
128'h06040513f00a15e310e91263470dd05c, /*  590 */
128'hd49b1ff4849b0024949bd408b17ff0ef, /*  591 */
128'h0793c45cc81c57fdee99e7e324810094, /*  592 */
128'h0654478308f91963478d00f402a3f800, /*  593 */
128'hd79b0107979b8fd90087979b06444703, /*  594 */
128'hf0ef8522001a859b06f71b6347054107, /*  595 */
128'h02a32324470323344783e13d2501ce5f, /*  596 */
128'hd79b776d0107979b8fd90087979b0004, /*  597 */
128'hf0ef0344051304f71263a55707134107, /*  598 */
128'h02f51763252787932501416157b7a99f, /*  599 */
128'h87932501614177b7a83ff0ef21840513, /*  600 */
128'hc808a6dff0ef21c4051300f51c632727, /*  601 */
128'hd78300009797c448a63ff0ef22040513, /*  602 */
128'h7cf719230000971793c117c227857e07, /*  603 */
128'hb351478100042a230124002300f41323, /*  604 */
128'h0513b5b90005099ba33ff0ef05840513, /*  605 */
128'hd41c9fb5e00a05e3b545a25ff0ef0544, /*  606 */
128'h87bb478db7010014949b00f915634789, /*  607 */
128'he8221101bdc59cbd0017d79b88850297, /*  608 */
128'h4703ed692501bffff0ef842ae426ec06, /*  609 */
128'h1b634785005447030cf71063478d0004, /*  610 */
128'hf0ef8526458120000613034404930af7, /*  611 */
128'h09a3faa0079322f4092305500793a01f, /*  612 */
128'h079302f40aa302f40a230520079322f4, /*  613 */
128'h04100713481c20f40da302f40b230610, /*  614 */
128'h0107571b0107971b20e40d2302e40ba3, /*  615 */
128'h0107d71b20e40ea320f40e230087571b, /*  616 */
128'h501020e40f23445c20f40fa30187d79b, /*  617 */
128'h001445030087571b0107571b0107971b, /*  618 */
128'hd71b260522e400a322f4002307200693, /*  619 */
128'h012320d40ca320d40c230187d79b0107, /*  620 */
128'h63d050ef85a64685d81022f401a322e4, /*  621 */
128'h631050ef4581460100144503000402a3, /*  622 */
128'h8082610564a2644260e200a035332501, /*  623 */
128'h0025458300f6f96337f9ffe5869b4d1c, /*  624 */
128'h47858082450180829d2d02d585bb5548, /*  625 */
128'hec26f022f406e84a71794d180eb7f763, /*  626 */
128'h842e46890005470302e5f963892ae44e, /*  627 */
128'hd49b00f71e6308d70e63468d06d70c63, /*  628 */
128'hac7ff0ef9dbd0094d59b9cad515c0015, /*  629 */
128'h69a2694264e2740270a257fdc9112501, /*  630 */
128'hd59b0014899b0249278380826145853e, /*  631 */
128'h0344c483854a9dbd94ca1ff4f4930099, /*  632 */
128'h4783994e1ff9f993f5792501a93ff0ef, /*  633 */
128'hbf658391c0198fc50087979b88050349, /*  634 */
128'h9dbd0085d59b515cbf458fe9157d6505, /*  635 */
128'h1fe474130014141bfd592501a63ff0ef, /*  636 */
128'h8fc90087979b03494503035947839922, /*  637 */
128'h2501a39ff0ef9dbd0075d59b515cb759, /*  638 */
128'h954a034505131fc575130024151bf935, /*  639 */
128'h4785b76517fd2501100007b7807ff0ef, /*  640 */
128'hf426fc06f04a4540f82271398082853e, /*  641 */
128'h1c63892a478500b51523e456e852ec4e, /*  642 */
128'h6a4269e2790274a2744270e2450900f4, /*  643 */
128'h84aefee474e34f98611c808261216aa2, /*  644 */
128'heb15579800e69463470d0007c683e021, /*  645 */
128'hd171008928235788fce4f7e30087d703, /*  646 */
128'h8793049688bd000937839d3d0044d79b, /*  647 */
128'hb75d450100993c2300a92a2394be0347, /*  648 */
128'h35034a8509925a7d843a0027c9838722, /*  649 */
128'hbf752501e59ff0ef0134f66385a20009, /*  650 */
128'hf68afbe301440c630005041be6fff0ef, /*  651 */
128'hbfc1413484bbf6f476e34f9c00093783, /*  652 */
128'hec06e426e822110100a55583b78d4505, /*  653 */
128'h6008484ce4950005049bf33ff0ef842a, /*  654 */
128'h020006136c08ec990005049b933ff0ef, /*  655 */
128'h601c00e7802357156c1cf3cff0ef4581, /*  656 */
128'h610564a28526644260e200e782234705, /*  657 */
128'hec4ef04af426f822fc06e85271398082, /*  658 */
128'hf063498984aa4d1c16ba75634a05e456, /*  659 */
128'h0ae78f63842e89324709000547830af5, /*  660 */
128'h515c0015da1b154794630ee78863470d, /*  661 */
128'h099b8b9ff0ef9dbd009a559b00ba0a3b, /*  662 */
128'h0ff97793001a0a9b8805060996630005, /*  663 */
128'h66850347c783014487b3cc191ffa7a13, /*  664 */
128'hf7938fd98ff50049179b00f7f71316c1, /*  665 */
128'h50dc00f48223478502fa0a239a260ff7, /*  666 */
128'h0005099b86bff0ef9dbd8526009ad59b, /*  667 */
128'h79130049591bc40d1ffafa9300099f63, /*  668 */
128'h70e200f482234785032a8a239aa60ff9, /*  669 */
128'h61216aa26a4269e2790274a2854e7442, /*  670 */
128'h79130089591b0347c783015487b38082, /*  671 */
128'h0085d59b515cb7e90127e9339bc100f9, /*  672 */
128'h141bfc0992e30005099b811ff0ef9dbd, /*  673 */
128'h0109191b03240a2394261fe474130014, /*  674 */
128'h0144822303240aa30089591b0109591b, /*  675 */
128'h099bfd8ff0ef9dbd0075d59b515cbf79, /*  676 */
128'h0a931fc474130024141bf80996e30005, /*  677 */
128'hf00006372501da0ff0ef85569aa60344, /*  678 */
128'h0107d79b94260109179b012569338d71, /*  679 */
128'h0109579b00fa80a30087d79b03240a23, /*  680 */
128'h4989b745012a81a300fa81230189591b, /*  681 */
128'he852f04af822fc06ec4ef4267139bf3d, /*  682 */
128'h04090a6300c52903e19d89ae84aae456, /*  683 */
128'h24054c9c5afd4a05844a04f977634d1c, /*  684 */
128'hc43ff0efa8214401052a606304f46363, /*  685 */
128'h00f41d6357fd0887f86347850005041b, /*  686 */
128'h6a4269e2790274a2744270e28522547d, /*  687 */
128'hb7d5faf47ee3894e4c9c808261216aa2, /*  688 */
128'h2501c05ff0ef852685a24409bf554905, /*  689 */
128'hb76dfb2411e305450863fd5507e3c901, /*  690 */
128'h2501de9ff0ef852685a2167d10000637, /*  691 */
128'hfae783e3577dc4c0489c02099063e905, /*  692 */
128'h00f482a30017e7930054c783c89c37fd, /*  693 */
128'hdd612501dbbff0ef852685ce8622bf49, /*  694 */
128'h5903f04a7139bfad4405f6f50fe34785, /*  695 */
128'hec4ef426030917932905f822fc0600a5, /*  696 */
128'h74a2744270e24511eb9993c1e456e852, /*  697 */
128'hd7ed495c808261216aa26a4269e27902, /*  698 */
128'h2785480c00099d63842a8a2e00f97993, /*  699 */
128'h75e30009071b00855783e18dc85c6108, /*  700 */
128'h97ce03478793012415230996601cfcf7, /*  701 */
128'h37fd00495a9b00254783bf5d4501ec1c, /*  702 */
128'h0005049bb27ff0effc0a9fe30157fab3, /*  703 */
128'h00f4946357fdbf4945090097e4634785, /*  704 */
128'hf60a0ee306f4e0634d1c6008b7614505, /*  705 */
128'h4785d4bd451d0005049be81ff0ef480c, /*  706 */
128'hdd8ff0ef6008fcf48de357fdfcf48be3, /*  707 */
128'h034505134581200006136008f5792501, /*  708 */
128'haa5ff0ef855285a600043a03beeff0ef, /*  709 */
128'h00faed630025478360084a0502aa2823, /*  710 */
128'hf0ef85a6c8046008d91c415787bb591c, /*  711 */
128'h2501d1cff0ef01450223b7b9c848a83f, /*  712 */
128'h7139b7e9db1c27855b1c2a856018f141, /*  713 */
128'he05ae456e852ec4ef04afc06f426f822, /*  714 */
128'h00e78663842e84aa02f007130005c783, /*  715 */
128'h47030004a62304050ce7906305c00713, /*  716 */
128'h05c00a9302f00a130ae7fc6347fd0004, /*  717 */
128'h80630d478263000447834b2102e00993, /*  718 */
128'hf0ef854a02000593462d0204b9030d57, /*  719 */
128'h4783013900230d37926300044783b40f, /*  720 */
128'h478300f900a302e007930b3790630014, /*  721 */
128'h0793943a09479763470d1b378e630024, /*  722 */
128'h2501adbff0ef8526458100f905a30200, /*  723 */
128'he96d2501cdaff0ef608848cc10051063, /*  724 */
128'hef918ba100b74783c7e5000747836c98, /*  725 */
128'h4603078507050cb78d6300b78593709c, /*  726 */
128'hf0ef85264581fed608e3fff7c683fff7, /*  727 */
128'h85264581b791c55c4bdc611cbf75dfdf, /*  728 */
128'h74a2744270e20004bc232501a85ff0ef, /*  729 */
128'h0405808261216b026aa26a4269e27902, /*  730 */
128'he06302000693f7578be3bf954709bf1d, /*  731 */
128'h45a147014681b7ad02400793943a12f6, /*  732 */
128'he793a8dd0505a0d14865020003134781, /*  733 */
128'h268500e50023954a9101020695130027, /*  734 */
128'h15630e50069300094503c6ed4711a06d, /*  735 */
128'h0027979b0165966300d90023469500d5, /*  736 */
128'h671300b6946345850037f6930ff7f793, /*  737 */
128'h16020087671300d7946346918bb10107, /*  738 */
128'h4511bf654701bdfd00e905a394329201, /*  739 */
128'hf713f4e518e34711c50500b7c783709c, /*  740 */
128'h0004bc230004a623cb890207f7930047, /*  741 */
128'h8b91b73d4515fb0dbf154501e80703e3, /*  742 */
128'hc503609cdbe58bc100b5c7836c8cfbf5, /*  743 */
128'h979b05659a63bdb9c4c8af2ff0ef0007, /*  744 */
128'h0017061b873245ad46a10ff7f7930027, /*  745 */
128'h06e3f4e374e300074703972293011702, /*  746 */
128'h151b02b6f263fd370ae3f95704e3f947, /*  747 */
128'h05130000851700054c634185551b0187, /*  748 */
128'h4519f11710e300088663000548830c65, /*  749 */
128'h051beea87ae30ff57513fbf7051bbd6d, /*  750 */
128'h0017e7933701eea866e30ff57513f9f7, /*  751 */
128'he44ee84aec26f0227179bdf90ff77713, /*  752 */
128'h484c49bd0e500913451184aef406842a, /*  753 */
128'he1292501afaff0ef6008a0b1c90de199, /*  754 */
128'h03f7f79300b7c783c3210007c7036c1c, /*  755 */
128'h0017b79317e18bfd0337806303270263, /*  756 */
128'h69a2694264e2740270a2450100979a63, /*  757 */
128'hd9452501c13ff0ef8522458180826145, /*  758 */
128'he82245811101bfe54511b7cd00042a23, /*  759 */
128'h0493e50d250188fff0ef842ae426ec06, /*  760 */
128'h6c1ced092501a8cff0ef6008484c0e50, /*  761 */
128'hf0ef85224585cb9900978d630007c783, /*  762 */
128'h60e2451d00f513634791dd792501bcdf, /*  763 */
128'hec06e426e82211018082610564a26442, /*  764 */
128'h6008484ce49d0005049bfa9ff0ef842a, /*  765 */
128'h020006136c08e0850005049ba42ff0ef, /*  766 */
128'h82aff0ef462d6c08700c84cff0ef4581, /*  767 */
128'h64a28526644260e200e782234705601c, /*  768 */
128'h45098082450900b7ed63478580826105, /*  769 */
128'h808261456a0269a2694264e2740270a2, /*  770 */
128'he052e44ee84af406ec26f02271794d1c, /*  771 */
128'hfa634c1c59fd4a05fcf5fde384ae842a, /*  772 */
128'h14630005091bec8ff0ef852285a600f4, /*  773 */
128'h460103390763fb490ce3bf7545010009, /*  774 */
128'h8a63481cf15d25018afff0ef852285a6, /*  775 */
128'h02a30017e79300544783c81c27850137, /*  776 */
128'hec2a7139b7594505bf5d0009049b00f4, /*  777 */
128'h426383eff0eff42ee432e82efc061028, /*  778 */
128'h00a78733050ecc678793000097970405, /*  779 */
128'h0023c319676200070023c31966226318, /*  780 */
128'h00f618634785cb114501e39897aa0007, /*  781 */
128'h612170e22501a0eff0ef0828080c4601, /*  782 */
128'hfca6e122e506f8ca7175bfe5452d8082, /*  783 */
128'h14050d634925e42ee8daecd6f0d2f4ce, /*  784 */
128'hf0ef1028002c8a7984aa89b200053023, /*  785 */
128'h1028083c65a2140910630005091b9d6f, /*  786 */
128'h4519e011e11964062501b6dff0efe4be, /*  787 */
128'h16634791c54dc3e101f9fa1301c9f793, /*  788 */
128'he949008a6a132501e75ff0ef102800f5, /*  789 */
128'h0713046007937aa2cfcd008a77936406, /*  790 */
128'h07a30004072300f40ca300f408a30210, /*  791 */
128'h0c2300040ba300040b2300e408230004, /*  792 */
128'h0f2300040ea300040e23000405a300e4, /*  793 */
128'hfc9fe0ef85a2000ac50300040fa30004, /*  794 */
128'h0aa300040a2300040da300040d234785, /*  795 */
128'h85ce04098b6300fa82230005099b0004, /*  796 */
128'h7522e9112501e3fff0ef030aab038556, /*  797 */
128'hc90d250183aff0ef0135262385da39fd, /*  798 */
128'h0049f993e3d98bc500b44783a895892a, /*  799 */
128'hf71300b44783f565a0854921f60981e3, /*  800 */
128'he3ad8b85000984630029f993e72d0107, /*  801 */
128'ha78385a279a2020a6a13c399008a7793, /*  802 */
128'hc503000485a3d09c01448523f4800309, /*  803 */
128'hdbbfe0ef01c40513c8c8f33fe0ef0009, /*  804 */
128'hb0230004ae230004a623c8880069d783, /*  805 */
128'h794674e6854a640a60aa00f494230134, /*  806 */
128'hb7e54911808261496b466ae67a0679a6, /*  807 */
128'hfc86e4d6e8d2eccef8a27119b7d5491d, /*  808 */
128'hec6ef06af466f862fc5ee0daf0caf4a6, /*  809 */
128'he91fe0ef8ab6e4328a2e842a0006a023, /*  810 */
128'hc39d662200b44783000998630005099b, /*  811 */
128'h69e6790674a6854e744670e60007899b, /*  812 */
128'h6de27d027ca27c427be26b066aa66a46, /*  813 */
128'h2903160789638b8500a4478380826109, /*  814 */
128'h091b00f67463893e40f907bb445c0104, /*  815 */
128'hfa090ce35c7d03040b1320000b930006, /*  816 */
128'h00975c9b6008120790631ff777934458, /*  817 */
128'h99630ffcfc930197fcb337fd00254783, /*  818 */
128'h05a3478900a7ec6347854848eb11020c, /*  819 */
128'hb7e52501bd6ff0ef4c0cb741498900f4, /*  820 */
128'hcc08b7a5498500f405a3478501851763, /*  821 */
128'hd5792501b98ff0ef856e4c0c00043d83, /*  822 */
128'h0007849b00a6073b0099579b000c861b, /*  823 */
128'h84bb00f6f4639fb1002dc683c4b58d3a, /*  824 */
128'h14a050ef85d2863a86a6001dc5034196, /*  825 */
128'h4c48c3850407f79300a44783f94d2501, /*  826 */
128'h910115020097951b0097fc6341a507bb, /*  827 */
128'h0094949bc5ffe0ef955285da20000613, /*  828 */
128'h9fa54099093b445c9a3e938102049793, /*  829 */
128'h4c50b70500faa0239fa5000aa783c45c, /*  830 */
128'hc503c38d0407f79300a4478304e60163, /*  831 */
128'hf1392501110050efe43a85da4685001d, /*  832 */
128'h601c00f40523fbf7f793672200a44783, /*  833 */
128'h25010bc050ef85da0017c503863a4685, /*  834 */
128'h1ff5f5930009049b444c01a42e23f115, /*  835 */
128'h030585930007849b0127f46340bb87bb, /*  836 */
128'hb59d499dbf9dbd1fe0ef855295a28626, /*  837 */
128'heca6f486fc56e0d2e4cee8caf0a27159, /*  838 */
128'h0006a023e46ee86aec66f062f45ef85a, /*  839 */
128'h0005099bcb5fe0ef8ab689328a2e842a, /*  840 */
128'h70a60007899bc39d00b4478300099763, /*  841 */
128'h7b427ae26a0669a6694664e6854e7406, /*  842 */
128'h4783808261656da26d426ce27c027ba2, /*  843 */
128'h6c630127873b445c18078f638b8900a4, /*  844 */
128'h046344585c7d03040b1320000b9304f7, /*  845 */
128'h00975c9b6008140793631ff777930409, /*  846 */
128'h9a630ffcfc930197fcb337fd00254783, /*  847 */
128'h02e798634705cb914581485cef01040c, /*  848 */
128'hd86ff0ef4c0cb759498900f405a34789, /*  849 */
128'h478312f76a634818445cf3fd0005079b, /*  850 */
128'h01879763b79500f405230207e79300a4, /*  851 */
128'he311cc1c4858bf99498500f405a34785, /*  852 */
128'h4c50601cc38d0407f79300a44783c85c, /*  853 */
128'hf96925017b1040ef85da0017c5034685, /*  854 */
128'h00043d8300f40523fbf7f79300a44783, /*  855 */
128'h000c869bd159250197cff0ef856e4c0c, /*  856 */
128'hc4b58d320007849b00a6863b0099579b, /*  857 */
128'hc503419704bb00f774639fb5002dc703, /*  858 */
128'h4c4cf1512501763040ef85d286a6001d, /*  859 */
128'h918115820097959b0297f26341a587bb, /*  860 */
128'h00a44783a4ffe0ef855a95d220000613, /*  861 */
128'h020497930094949b00f40523fbf7f793, /*  862 */
128'ha783c45c9fa54099093b445c9a3e9381, /*  863 */
128'h00c78e634c5cbdd100faa0239fa5000a, /*  864 */
128'h85da4685001dc50300e7fa63445c4818, /*  865 */
128'h049b444801a42e23fd0925016c7040ef, /*  866 */
128'h849b0127f46340ab87bb1ff575130009, /*  867 */
128'h9dbfe0ef952285d28626030505130007, /*  868 */
128'hc81cbf4100f405230407e79300a44783, /*  869 */
128'he0ef842ae406e0221141bd2d499db5f9, /*  870 */
128'hcf690207f71300a44783e1752501acff, /*  871 */
128'h0017c50346854c50601cc3950407f793, /*  872 */
128'h00a44783ed552501685040ef03040593, /*  873 */
128'hb77fe0ef6008500c00f40523fbf7f793, /*  874 */
128'h85a30207671300b7c703741ce15d2501, /*  875 */
128'h0086d69b0106d69b0107169b481800e7, /*  876 */
128'h0187571b0107569b00d78ea300e78e23, /*  877 */
128'h8ba300078b23485800e78fa300d78f23, /*  878 */
128'h27010107571b0107169b00e78d230007, /*  879 */
128'h0087571b0107571b0107171b00e78a23, /*  880 */
128'h00e78c23021007130106d69b00e78aa3, /*  881 */
128'h00e78ca300d78da3046007130086d69b, /*  882 */
128'hf793600800a44783000789a300078923, /*  883 */
128'h60a2640200f50223478500f40523fdf7, /*  884 */
128'h80820141640260a24505ebbfe06f0141, /*  885 */
128'he9012501effff0ef842ae406e0221141, /*  886 */
128'h60a200043023e11925019cbfe0ef8522, /*  887 */
128'he0efec060028e42a1101808201416402, /*  888 */
128'h45015ea789230000879700054a6395bf, /*  889 */
128'h4601e42a7159bfe5452d8082610560e2, /*  890 */
128'h041bb3bfe0efeca6f486f0a21028002c, /*  891 */
128'hcd2ff0efe4be1028083c65a2ec190005, /*  892 */
128'hcbd8575277a2e9916586e41d0005041b, /*  893 */
128'h00b5c7838082616564e6740670a68522, /*  894 */
128'hc8c897bfe0ef0004c50374a2cb998bc1, /*  895 */
128'hfca67175bfd94415fcf41ee34791b7c5, /*  896 */
128'h00050023f0d2f4cef8cae122e506e42a, /*  897 */
128'he5292501acdfe0ef1828002c460184ae, /*  898 */
128'h02f009934bdc597d842677e2ecbe081c, /*  899 */
128'h8717e50567a24501040a12634a16c2be, /*  900 */
128'h071300e780230307071b53a747030000, /*  901 */
128'h812302f007130e94186300e780a303a0, /*  902 */
128'h794674e6640a60aa00078023078d00e7, /*  903 */
128'hf89fe0ef18284585808261497a0679a6, /*  904 */
128'hf5552501e6eff0ef18284581fd452501, /*  905 */
128'h4581c2aa8cdfe0ef0007c50365c677e2, /*  906 */
128'hf0ef18284581f9492501f63fe0ef1828, /*  907 */
128'he0ef0007c50365c677e2e1052501e48f, /*  908 */
128'ha9eff0ef1828458101450e6325018a7f, /*  909 */
128'hb7594509f8e516e367a24711dd612501, /*  910 */
128'h9301020797134781f5cfe0ef1828100c, /*  911 */
128'h62630037871beb05fc97470397361094, /*  912 */
128'h961300e586bb40f405bbfff7871b04e4, /*  913 */
128'hfff7c79301271a6396b2920166a20206, /*  914 */
128'h02071613b7c12785b7319c3d01368023, /*  915 */
128'h00c68023377dfc964603962a10889201, /*  916 */
128'h92810204169367220789bddd4545b7e9, /*  917 */
128'h65e3fee78fa324050785000747039736, /*  918 */
128'hec4efc06f04af426f8227139b709fe94, /*  919 */
128'h0005091bfb4fe0ef84ae842ae456e852, /*  920 */
128'h70e20007891bcf8900b4478300091763, /*  921 */
128'h61216aa26a4269e2790274a2854a7442, /*  922 */
128'he3918b8900a447830097776348188082, /*  923 */
128'h78e34818445ce4bd00042623445884ba, /*  924 */
128'h00f405230207e79300a44783c81cfcf7, /*  925 */
128'h0ee34c50d3e51ff7f793445c4481bf7d, /*  926 */
128'hc3850407f7930304099300a44783fc96, /*  927 */
128'h250130f040ef0017c50385ce4685601c, /*  928 */
128'h601c00f40523fbf7f79300a44783ed51, /*  929 */
128'h25012bd040ef85ce0017c50386264685, /*  930 */
128'h0097999b002547836008bf59cc44ed35, /*  931 */
128'h0337563b0336d6bbfff4869b377dc729, /*  932 */
128'hc45c27814c0c8ff9413007bb02c6ed63, /*  933 */
128'h9fa5445c0499ea634a855a7dd1c19c9d, /*  934 */
128'h2501c87fe0ef6008d7b51ff4f793c45c, /*  935 */
128'hf0efe595484cbfb19ca90094d49bcd11, /*  936 */
128'h05a3478900f5976347850005059b814f, /*  937 */
128'h05a3478500f5976357fdbded490900f4, /*  938 */
128'h00a44783b765cc0cc84cb5ed490500f4, /*  939 */
128'he5990005059bfddfe0efcb818b896008, /*  940 */
128'hfd4588e30005059bc4bfe0efbf6984ce, /*  941 */
128'hcc0c445cfaf5fae34f9c601cfabafee3, /*  942 */
128'hfc067139b7bdc45c013787bb413484bb, /*  943 */
128'he0ef0828002c4601842ac52de42ef822, /*  944 */
128'h101ce01c852265a267e2e1152501fe6f, /*  945 */
128'hc783cd996c0ce529250197cff0eff01c, /*  946 */
128'h67e2a02d000430234515e7898bc100b5, /*  947 */
128'h8522458167e2c448e30fe0ef0007c503, /*  948 */
128'h47912501cbdfe0ef00f414230067d783, /*  949 */
128'h452580826121744270e2f971fcf50be3, /*  950 */
128'he406e0221141b7c1fcf501e34791bfdd, /*  951 */
128'h60a200043023e1192501dbafe0ef842a, /*  952 */
128'hf406e84aec26f0227179808201416402, /*  953 */
128'h1f63e8890005049bd98fe0ef892e842a, /*  954 */
128'h70a20005049bc5ffe0ef852245810009, /*  955 */
128'h022430238082614564e2694285267402, /*  956 */
128'h02f5136347912501b32ff0ef85224581, /*  957 */
128'h85224581c68fe0ef852285ca00042a23, /*  958 */
128'h00042a2300f5166347912501f8bfe0ef, /*  959 */
128'h84aee42aeca67159bf6584aad16dbf7d, /*  960 */
128'h041bedafe0eff486f0a21028002c4601, /*  961 */
128'h872ff0efe4be1028083c65a2e00d0005, /*  962 */
128'h102885a6c489cf816786e8010005041b, /*  963 */
128'h8082616564e6740670a68522c10fe0ef, /*  964 */
128'h8b2ee42af85a8432f0a27159bfcd4419, /*  965 */
128'he4cee8caeca6f486e0d28522002c4601, /*  966 */
128'h00050a1be7cfe0efec66f062f45efc56, /*  967 */
128'hffec871b481c01842c836000000a1c63, /*  968 */
128'h64e68552740670a600fb202302f76263, /*  969 */
128'h6ce27c027ba27b427ae26a0669a66946, /*  970 */
128'h490902fb9f63478500044b8380826165, /*  971 */
128'h2501a55fe0ef852285ca4a8559fd4481, /*  972 */
128'h29054c1c2485e1110955086309350863, /*  973 */
128'h02a30017e793c80400544783fef963e3, /*  974 */
128'h490110000ab7504cb74d009b202300f4, /*  975 */
128'h899b852200099e631afd4c0944814981, /*  976 */
128'h0344091385cee9212501d10fe0ef0015, /*  977 */
128'h0009470300194783038b916320000993, /*  978 */
128'h3cfd39f909092485e3918fd90087979b, /*  979 */
128'h2501abcfe0efe02e854ab745fc0c94e3, /*  980 */
128'hb7c539f109112485e111658201557533, /*  981 */
128'he8221101bfad8a2abfbd4a09b7494a05, /*  982 */
128'h0005049bbc4fe0ef842ae04aec06e426, /*  983 */
128'h644260e20007849bcb9100b44783e491, /*  984 */
128'hf71300a447838082610564a269028526, /*  985 */
128'h0207e793fed772e348144458cf390027, /*  986 */
128'ha58ff0ef484cef01600800f40523c818, /*  987 */
128'hbf7d84aa00a405a3c53900042a232501, /*  988 */
128'h02f9146357fd0005091b94dfe0ef4c0c, /*  989 */
128'hb37fe0ef167d100006374c0cb7dd4505, /*  990 */
128'hb7e12501a1cff0ef85ca6008f9792501, /*  991 */
128'h4d1c6008fcf900e345094785b769449d, /*  992 */
128'h601cdba50407f79300a44783fcf96ae3, /*  993 */
128'h6ec040ef030405930017c50346854c50, /*  994 */
128'h00f40523fbf7f79300a44783f55d2501, /*  995 */
128'he122e5061008002c4605e42a7175b7b1, /*  996 */
128'h081c65a2e9052501ca0fe0eff8cafca6, /*  997 */
128'h45196786e1052501e3bfe0efe0be1008, /*  998 */
128'hc483c59975e2eb890207f79300b7c783, /*  999 */
128'h74e6640a60aa451dcb810014f79300b5, /* 1000 */
128'had8fe0ef000945037902808261497946, /* 1001 */
128'h8de301492783c89d88c1cc0d0005041b, /* 1002 */
128'h458996cfe0ef00a8100c02800613fc87, /* 1003 */
128'h00a84581f1612501951fe0efcaa200a8, /* 1004 */
128'h1008faf518e34791d94d2501836ff0ef, /* 1005 */
128'hf20fe0ef7502e411f15525019f5fe0ef, /* 1006 */
128'hd575250191cff0ef85a27502bf612501, /* 1007 */
128'hf506f1221028002c4605e42a7171b769, /* 1008 */
128'hf0e2f4def8dafcd6e152e54ee94aed26, /* 1009 */
128'h1c0414630005041bbd0fe0efe8eaece6, /* 1010 */
128'h0005041bd67fe0efe4be1028083c65a2, /* 1011 */
128'hc783441967a61af4176347911c040963, /* 1012 */
128'he0ef4581752218079f630207f79300b7, /* 1013 */
128'h0f6344094785180902630005091bb45f, /* 1014 */
128'ha98fe0ef752216f90b63440557fd16f9, /* 1015 */
128'h0109549b85ca7422160414630005041b, /* 1016 */
128'h45812000061303440a13f6efe0ef8522, /* 1017 */
128'h02000593462d898fe0ef855200050c1b, /* 1018 */
128'h199b0ff4fb1347c1248188cfe0ef8552, /* 1019 */
128'h07930109d99b02f40fa30104949b0109, /* 1020 */
128'h7a9304f4062302e00b930104d49b0210, /* 1021 */
128'h06a30084d49b0089d99b046007930ff9, /* 1022 */
128'h05a30404052303740a230200061304f4, /* 1023 */
128'h04a305640423053407a3055407230404, /* 1024 */
128'h0aa3772280efe0ef0544051385d20494, /* 1025 */
128'h571400d6166357d200074603468d0574, /* 1026 */
128'hd79b0107969b06f40723478100f69363, /* 1027 */
128'h0106d69b0107979b06f4042327810107, /* 1028 */
128'h06d407a30087d79b0086d69b0107d79b, /* 1029 */
128'h1028040b99634c8500274b8306f404a3, /* 1030 */
128'h752247416786e8350005041bf59fe0ef, /* 1031 */
128'h0460071300e78c230210071300e785a3, /* 1032 */
128'h01578d2300e78ca300078ba300078b23, /* 1033 */
128'h0223478500978aa301678a2301378da3, /* 1034 */
128'h0d1b7522a82d0005041bd5afe0ef00f5, /* 1035 */
128'h041b8dcfe0ef0195022303852823001c, /* 1036 */
128'hd0ef3bfd8552458120000613ec090005, /* 1037 */
128'h85ca7522441db7498c6a0ffbfb93f61f, /* 1038 */
128'h69aa694a64ea740a70aa8522f25fe0ef, /* 1039 */
128'h614d6d466ce67c067ba67b467ae66a0a, /* 1040 */
128'h84aee42aeca6f0a27159b7c544218082, /* 1041 */
128'h25019cafe0eff48610284605002c8432, /* 1042 */
128'h2501b65fe0efe4be1028083c65a2e131, /* 1043 */
128'he39d0207f79300b7c783451967a6e915, /* 1044 */
128'h74138c658cbd752200b74783c30d6706, /* 1045 */
128'he0ef00f502234785008705a38c3d0274, /* 1046 */
128'h71718082616564e6740670a62501c9ef, /* 1047 */
128'hed26f122f5060088002c4605e02ee42a, /* 1048 */
128'h65a26786120796630005079b964fe0ef, /* 1049 */
128'h0005079baf7fe0eff0be083cf4be0088, /* 1050 */
128'h02077713479900b7c703778610079a63, /* 1051 */
128'h05ad46550e058e63479165e610071263, /* 1052 */
128'hd0ef10a8008c02800613e55fd0ef1028, /* 1053 */
128'h65820c054d6347adf05fd0ef850ae49f, /* 1054 */
128'h93634711cbf90005079baadfe0ef10a8, /* 1055 */
128'h648aefc50005079bdc5fe0ef10a80ce7, /* 1056 */
128'h4783e0dfd0ef00d4851302a10593464d, /* 1057 */
128'h0223478500f485a30207e79364060281, /* 1058 */
128'h086357d64736cbbd8bc100b4c78300f4, /* 1059 */
128'h0005059bf2dfd0ef85a60004450306f7, /* 1060 */
128'h8522c5a547890005059bcaefe0ef8522, /* 1061 */
128'h02e007936706efb10005079bfc3fd0ef, /* 1062 */
128'h07230107969b57d602f69d6305574683, /* 1063 */
128'h0107979b06f7042327810107d79b06f7, /* 1064 */
128'h0086d69b0106d69b0087d79b0107d79b, /* 1065 */
128'h008800f7022306d707a3478506f704a3, /* 1066 */
128'hb50fe0ef6506e7910005079be24fe0ef, /* 1067 */
128'h8082614d853e64ea740a70aa0005079b, /* 1068 */
128'h002c4605842ee42ae8a2711dbfcd47a1, /* 1069 */
128'h083c65a2e9292501810fe0efec861028, /* 1070 */
128'h451967a6e12925019abfe0efe4be1028, /* 1071 */
128'h5703cb856786eb950207f79300b7c783, /* 1072 */
128'h00e78ba30087571b00e78b2375220064, /* 1073 */
128'h00e78ca30087571b00e78c2300445703, /* 1074 */
128'h644660e62501ad6fe0ef00f502234785, /* 1075 */
128'h893284aee42ae0cae4a6711d80826125, /* 1076 */
128'h041bf9bfd0efec86e8a208284601002c, /* 1077 */
128'hca8fe0efd20208284581c4b9e0510005, /* 1078 */
128'he93d2501b8ffe0ef08284585e5592501, /* 1079 */
128'h46ad00b48713ca1fd0ef8526462d75c2, /* 1080 */
128'h869bfff6879bce890007002302000613, /* 1081 */
128'h83e3177d0007c78397a6938117820007, /* 1082 */
128'h041be69fd0ef510c656202090a63fec7, /* 1083 */
128'h0005468304300793470d6562e0150005, /* 1084 */
128'hd0ef953e034787930270079300e68463, /* 1085 */
128'h690664a6644660e6852200a92023c29f, /* 1086 */
128'hbf550004802300f51563479180826125, /* 1087 */
128'he8a21028002c4605e42a711db7d5842a, /* 1088 */
128'h0c2366a2ec550005041bee3fd0efec86, /* 1089 */
128'h0007c78397b693810206179346010001, /* 1090 */
128'he0efda0210284581ea2902000593eba1, /* 1091 */
128'habbfe0ef10284585e8410005041bbd6f, /* 1092 */
128'h082c462dc3dd650601814783e1792501, /* 1093 */
128'h071300e78c23021007136786bc7fd0ef, /* 1094 */
128'ha06100e78ca300078ba300078b230460, /* 1095 */
128'h02079713fff6079bbf45863eb74d2605, /* 1096 */
128'h4781082cfeb706e30007470397369301, /* 1097 */
128'h27850006c70348b107f00e9343658e2e, /* 1098 */
128'h1742370100a36c6391411542f9f7051b, /* 1099 */
128'ha82100070f1bade50513000075179341, /* 1100 */
128'h80826125644660e68522441900eef863, /* 1101 */
128'h1be306080563000548030505bfcdf36d, /* 1102 */
128'ha885078500c6802300fe06b3b7cdffe8, /* 1103 */
128'he0ef00f502234785752200f500235795, /* 1104 */
128'h478302f51b634791b7c10005041b8fef, /* 1105 */
128'hf4450005041ba55fe0ef1028dbd50181, /* 1106 */
128'h462d6506b07fd0ef4581020006136506, /* 1107 */
128'hbf1900e785a347216786ae5fd0ef082c, /* 1108 */
128'h0585068500e58023f91780e3b751842a, /* 1109 */
128'h869b02000613472993811782f4c7e5e3, /* 1110 */
128'h1de30e50079301814703f8d771e30007, /* 1111 */
128'h0585230305452e0305052e83bf89eaf7, /* 1112 */
128'h02938f2ae44ae826ec22110105c52883, /* 1113 */
128'h8f9300005f97887687f2869a86460405, /* 1114 */
128'h000fa38300b647338dfd00c6c5b3656f, /* 1115 */
128'h9db9007585bb0fc1008fa403000f2583, /* 1116 */
128'h0078159b0105883b004f2703ff4fa383, /* 1117 */
128'h00f805bb0077073b0105e8330198581b, /* 1118 */
128'h9e39008f23838e358e6d00f6c6339f31, /* 1119 */
128'h873b008383bb8e590146561b00c6171b, /* 1120 */
128'h00cf24038ef900b7c6b300d383bb00c5, /* 1121 */
128'he6b30116969b00f6d39b007686bb8ebd, /* 1122 */
128'h0007061b00d703bbffcfa4039fa100d3, /* 1123 */
128'h00a7579b9f3d8f2d9fa1007777338f2d, /* 1124 */
128'h0003869b0005881b0f418f5d0167171b, /* 1125 */
128'h6985859300005597f45f17e300e387bb, /* 1126 */
128'h69828293000052975d0f8f9300005f97, /* 1127 */
128'h000faf0301e6c73300cf7f3300d7cf33, /* 1128 */
128'h0005c70300ef0f3b0025c4030015c383, /* 1129 */
128'h0f3b942a040a4318972a070a93aa038a, /* 1130 */
128'h9e3900581f1b010f083b004fa70300ef, /* 1131 */
128'h00f80f3b010f68330003a70301b8581b, /* 1132 */
128'h008fa7039e398e3d8e7501e7c6339f31, /* 1133 */
128'h00c3e63340189eb90176561b0096139b, /* 1134 */
128'hc4838efd007f46b305919f3500cf03bb, /* 1135 */
128'h048affcfa7039eb90fc101e6c6b3fff5, /* 1136 */
128'h8ec140980126d69b9fb900e6941b94aa, /* 1137 */
128'h473301e777330083c7339fb900d3843b, /* 1138 */
128'h081b8f5d0147171b00c7579b9f3d0077, /* 1139 */
128'h99e300e407bb0004069b0003861b000f, /* 1140 */
128'h000053978ffa5aef0f1300005f17f255, /* 1141 */
128'h00d7c2b30003a703010fc40352438393, /* 1142 */
128'h011fc4839f25400000c2c4b3942a040a, /* 1143 */
128'h083b40809e2194aa048a0043a4039f21, /* 1144 */
128'h683301c8581b0048171b012fc4830107, /* 1145 */
128'hc2b3048a00f8073b0083a4039e210107, /* 1146 */
128'h00b6129b408000c2863b9ea194aa00e2, /* 1147 */
128'h02bb03c100c2e6330156561b013fc903, /* 1148 */
128'h0056c6b300e7c6b3ffc3a4839c3500c7, /* 1149 */
128'h0106d69b9fa50106941b992a9ea1090a, /* 1150 */
128'h47330007081b00d2843b8ec100092483, /* 1151 */
128'h0177171b0097579b9f3d8f219fa50057, /* 1152 */
128'h00e407bb0004069b0002861b0f918f5d, /* 1153 */
128'hfff6471349c2829300005297f5f592e3, /* 1154 */
128'h4403021f43830002a70300d745b38f5d, /* 1155 */
128'h95aa058a93aa038a020f45839f2d022f, /* 1156 */
128'h0107083b0042a5839f2d942a040a418c, /* 1157 */
128'h683301a8581b0003a5839e2d0068171b, /* 1158 */
128'h8e3d8e59fff6c6139db100f8073b0107, /* 1159 */
128'h9ead0166561b00a6139b0082a5839e2d, /* 1160 */
128'h023f44839ead00c703bb00c3e633400c, /* 1161 */
128'hffc2a4038db902c10075e5b3fff7c593, /* 1162 */
128'h8dd50115d59b94aa00f5969b048a9db5, /* 1163 */
128'hfff747130007081b00b385bb40809fa1, /* 1164 */
128'h171b00b7579b9f3d007747339fa18f4d, /* 1165 */
128'h87bb0005869b0003861b0f118f5d0157, /* 1166 */
128'h00fe07bb010e883b6462f3ef9de300e5, /* 1167 */
128'hcd34c97c0505282300c8863b00d306bb, /* 1168 */
128'he0a2715d653c80826105692264c2cd70, /* 1169 */
128'hec56f052e486e45ee85af44ef84afc26, /* 1170 */
128'h0b13e53c893289ae84aa97b203f7f413, /* 1171 */
128'h178200078a1b408b07bb04000b930400, /* 1172 */
128'hda93020a1a9300090a1b00f974639381, /* 1173 */
128'h20ef0144043b86560084853385ce020a, /* 1174 */
128'h852660bc0174176399d6415909334810, /* 1175 */
128'h79a2794274e2640660a6b7c997824401, /* 1176 */
128'h7179653c808261616ba26b426ae27a02, /* 1177 */
128'he84af406e44eec26842a03f7f793f022, /* 1178 */
128'h099300e7802397a2f800071300178513, /* 1179 */
128'h920116020006091b40a9863b449d0400, /* 1180 */
128'h078e643c0124f5633c9020ef95224581, /* 1181 */
128'h70a2fd24fde3450197828522603cfc1c, /* 1182 */
128'h000077978082614569a2694264e27402, /* 1183 */
128'h00007797e93c04053423639c14478793, /* 1184 */
128'hb6c7879300000797ed3c639c13c78793, /* 1185 */
128'hec06850a46410505059311018082e13c, /* 1186 */
128'h659735a686930000769747013bf020ef, /* 1187 */
128'h0007c78300e107b34541572585930000, /* 1188 */
128'h000646038bbd962e0047d61307050689, /* 1189 */
128'h1de3fef68fa3fec68f230007c78397ae, /* 1190 */
128'h8082610531c505130000751760e2fca7, /* 1191 */
128'hf71ff0efe42ee5060808842ae1227175, /* 1192 */
128'hf01ff0ef0808e85ff0ef080885a26622, /* 1193 */
128'h595880826149640a60aaf83ff0ef0808, /* 1194 */
128'h071300d71763469100d70d63711c46a1, /* 1195 */
128'h556dbfe50007ac2380824501cf980200, /* 1196 */
128'h842a420007b7ec06e426e82211018082, /* 1197 */
128'h061324a686930000569702f5026384ae, /* 1198 */
128'h0513000065174d658593000065970880, /* 1199 */
128'h610564a2644260e2fc2419b030ef4e65, /* 1200 */
128'h420007b7ec06e4266100e82211018082, /* 1201 */
128'h0613222686930000569702f4026384ae, /* 1202 */
128'h051300006517496585930000659702f0, /* 1203 */
128'h610564a2644260e2e00415b030ef4a65, /* 1204 */
128'h420007b7ec06e4266100e82211018082, /* 1205 */
128'h06131f2686930000569702f4026384ae, /* 1206 */
128'h05130000651745658593000065970360, /* 1207 */
128'h610564a2644260e2e40411b030ef4665, /* 1208 */
128'h420007b7ec06e8226104e42611018082, /* 1209 */
128'h061309a686930000769702f48263842e, /* 1210 */
128'h051300006517416585930000659703e0, /* 1211 */
128'h644260e2e880900114020db030ef4265, /* 1212 */
128'hec06e8226104e42611018082610564a2, /* 1213 */
128'h86930000769702f48263842e420007b7, /* 1214 */
128'h65173d258593000065970450061304e6, /* 1215 */
128'hec8090011402097030ef3e2505130000, /* 1216 */
128'h6100e82211018082610564a2644260e2, /* 1217 */
128'h569702f4026384ae420007b7ec06e426, /* 1218 */
128'h85930000659704c0061313a686930000, /* 1219 */
128'hf004053030ef39e505130000651738e5, /* 1220 */
128'h6100e82211018082610564a2644260e2, /* 1221 */
128'h569702f4026384ae420007b7ec06e426, /* 1222 */
128'h8593000065970530061310a686930000, /* 1223 */
128'hf404013030ef35e505130000651734e5, /* 1224 */
128'h3983ec4e71398082610564a2644260e2, /* 1225 */
128'h84ae420007b7fc06f04af426f8220005, /* 1226 */
128'h0d0686930000569702f9846384368932, /* 1227 */
128'h00006517304585930000659705a00613, /* 1228 */
128'h0014159b67227c6030efe43a31450513, /* 1229 */
128'h949b8dd9004979130029191b8b058989, /* 1230 */
128'hb8238dc5744270e288a10125e5b30034, /* 1231 */
128'he02211418082612169e2790274a202b9, /* 1232 */
128'hf0efe406458185224605468147057100, /* 1233 */
128'h468547058522f35ff0ef45818522f7df, /* 1234 */
128'hd97ff0ef45816008f67ff0ef45814605, /* 1235 */
128'he022e4061141808201414501640260a2, /* 1236 */
128'h45810405302302053c23460546814705, /* 1237 */
128'h8522ef1ff0ef45818522f39ff0ef842a, /* 1238 */
128'h64026008f23ff0ef4605468547054581, /* 1239 */
128'h6104e4261101d4dff06f0141458160a2, /* 1240 */
128'h569702f48263842e420007b7ec06e822, /* 1241 */
128'h85930000659706100613ffa686930000, /* 1242 */
128'h14426e2030ef22e505130000651721e5, /* 1243 */
128'h11018082610564a2644260e2fc809041, /* 1244 */
128'h8263842e420007b7ec06e8226104e426, /* 1245 */
128'h659706800613fc6686930000569702f4, /* 1246 */
128'h30ef1ea50513000065171da585930000, /* 1247 */
128'h64a2644260e2e0a08c7d17fd678569e0, /* 1248 */
128'h07b7ec06e4266100e822110180826105, /* 1249 */
128'hf90686930000569702f4026384ae4200, /* 1250 */
128'h00006517194585930000659706f00613, /* 1251 */
128'h64a2644260e2e424658030ef1a450513, /* 1252 */
128'he426e82200053903e04a110180826105, /* 1253 */
128'h569702f9026384ae842a420007b7ec06, /* 1254 */
128'h85930000659707600613f5a686930000, /* 1255 */
128'h3c23612030ef15e505130000651714e5, /* 1256 */
128'h80826105690264a2644260e2c8440499, /* 1257 */
128'he0d2e4cef486e8caeca67100f0a27159, /* 1258 */
128'hd783020408a3ec66f062f45ef85afc56, /* 1259 */
128'h051345814611d01ce03084b2892e0005, /* 1260 */
128'hf0ef458560080e049c636ca020ef00c9, /* 1261 */
128'h9a6304043a03420007b700043983bf5f, /* 1262 */
128'h8b89c7090017f71344810049278316f9, /* 1263 */
128'h09638cdd03243c234c1c4485e391448d, /* 1264 */
128'h0144e493160786638b85008a2783000a, /* 1265 */
128'h4581d71ff0ef85224581460546814705, /* 1266 */
128'h00005c17852200892583be1ff0ef8522, /* 1267 */
128'h6a17852200095583c4fff0efed4c0c13, /* 1268 */
128'hf0ef852285a6c81ff0ef07aa0a130000, /* 1269 */
128'h460546854705cf5ff0ef85224581cbdf, /* 1270 */
128'h24058593000f45b7d27ff0ef85224581, /* 1271 */
128'hb583cd1ff0ef85224585e93ff0ef8522, /* 1272 */
128'hf0ef25810015e593009899b785220d89, /* 1273 */
128'h485c03aa8a9300006a9768198993eb7f, /* 1274 */
128'h7ae26a0669a6694664e6740670a6efe9, /* 1275 */
128'h44cc8082616545016ce27c027ba27b42, /* 1276 */
128'hdf3ff0ef8522488cdb7ff0efe0248522, /* 1277 */
128'h654100043883603cee079be38b85449c, /* 1278 */
128'h0e37431147014781458163900107e683, /* 1279 */
128'h00064803ec0689e36e89f005051300ff, /* 1280 */
128'h27810107e7b301e8183b070500371f1b, /* 1281 */
128'h971b0187d81bf2e50067036316fd0605, /* 1282 */
128'hd79b01c878330087981b010767330187, /* 1283 */
128'h170200be873b8fd98fe9010767330087, /* 1284 */
128'h470147812585e31c9746938183751782, /* 1285 */
128'h659714900613d766869300005697b765, /* 1286 */
128'h30eff6a5051300006517f5a585930000, /* 1287 */
128'h42000bb78b4ebd6100c4e493bd8541e0, /* 1288 */
128'h6517d5a5859300005597000b1d633b7d, /* 1289 */
128'h00043903b7116f6000eff5a505130000, /* 1290 */
128'h30ef855685d20f20061386e201790963, /* 1291 */
128'h8e6324818cfd4c81485c070934833de0, /* 1292 */
128'h7c1c00f76f630c893783020937031204, /* 1293 */
128'hb6fff0ef85224581cc5cf9200793c781, /* 1294 */
128'h2903c3950044f793b27ff0ef85224581, /* 1295 */
128'hf0ef85ca00896913ff39791385220144, /* 1296 */
128'h680000efefc505130000651785cad47f, /* 1297 */
128'hff397913852201442903c3950084f793, /* 1298 */
128'h0000651785cad1fff0ef85ca00496913, /* 1299 */
128'h3c83cfb50014f793658000efefc50513, /* 1300 */
128'h869300005697017c8c63038439030004, /* 1301 */
128'h7c1c332030ef855685d209c00613cc66, /* 1302 */
128'h0037f693470d02043c2300492783cba9, /* 1303 */
128'h480d468100c90793018c871308e69f63, /* 1304 */
128'h8763c3900086161bff87051363104591, /* 1305 */
128'h872a2685c3988f518361ff8737030106, /* 1306 */
128'h0027e793485ccbb5603cfeb690e30791, /* 1307 */
128'h6004cc9d4c858889c85c9bf9485cc85c, /* 1308 */
128'hc60686930000569701748c6304043903, /* 1309 */
128'h040430232b4030ef855685d20ca00613, /* 1310 */
128'hf0ef8522ef8d8b850089278300090963, /* 1311 */
128'hf0ef8522484cc85c9bf54c85485cb4df, /* 1312 */
128'h8b85bd95641020ef4505d80c8ee3c47f, /* 1313 */
128'hf0ef8522b77100f92623000cb783dbd9, /* 1314 */
128'h00093c830109648397a667a1bf41b1df, /* 1315 */
128'h46218566639c00878913fa978de394be, /* 1316 */
128'h5535b7dd87ca0ca139a020efe43e002c, /* 1317 */
128'he84aec26f02204800513717908b04163, /* 1318 */
128'h5551842a1a4030ef892e84b2e44ef406, /* 1319 */
128'h785010efbcc505130000551785a2cc1d, /* 1320 */
128'h00efdca5051300006517862285aa89aa, /* 1321 */
128'h01242423e01c420007b702098b634fe0, /* 1322 */
128'h70a24501c45c4789cb990024f793f404, /* 1323 */
128'h450188858082614569a2694264e27402, /* 1324 */
128'h557d18c030ef8522b7e5c45c4785d4fd, /* 1325 */
128'hf73ff06f42000537458146098082bff9, /* 1326 */
128'h711c808225016108953e050e420007b7, /* 1327 */
128'h02f40263420007b7e4066380e0221141, /* 1328 */
128'h0000659734c00613b686869300005697, /* 1329 */
128'h170030efcbc5051300006517cac58593, /* 1330 */
128'h80820141640260a2557de3914505703c, /* 1331 */
128'h4d3010efe42eec064501842ae8221101, /* 1332 */
128'h7940006f6105468560e26622644285a2, /* 1333 */
128'he44ee84aec26f022f406200005137179, /* 1334 */
128'hd20505130000651784aa0aa030efe052, /* 1335 */
128'h10ef450144b010ef0001b5031b2030ef, /* 1336 */
128'h051300006517681c206010ef842a4910, /* 1337 */
128'h0000651706f445833f8000ef638cd065, /* 1338 */
128'h051300006517546c3e8000efd0450513, /* 1339 */
128'h583c3d2000ef91c115c20085d59bd0e5, /* 1340 */
128'h0087d71bd04505130000651706c44583, /* 1341 */
128'h0ff7f7930ff777130187d61b0107d69b, /* 1342 */
128'h000065175c0c3a6000ef26010ff6f693, /* 1343 */
128'h859300006597545c398000efcf450513, /* 1344 */
128'h00006517c6c5859300006597c789c7e5, /* 1345 */
128'hcf05051300006517378000efce450513, /* 1346 */
128'hb0ef2f258593000065977448102030ef, /* 1347 */
128'hc486061300006617584c19c42783dbbf, /* 1348 */
128'h051300006517fa66061300006617e789, /* 1349 */
128'hed5ff0ef84264581852633a000efcce5, /* 1350 */
128'h899300006997ccea0a1300006a174481, /* 1351 */
128'h855285a6e78901f4f79320000913cce9, /* 1352 */
128'h00f5f6132485854e0004458330c000ef, /* 1353 */
128'h00006517fd249fe304052fa000ef8191, /* 1354 */
128'h694264e2740270a22e8000ef27c50513, /* 1355 */
128'hb7830103b7038082614545016a0269a2, /* 1356 */
128'h93811782278540f707b30003b6830083, /* 1357 */
128'h00a7002300f3b8230017079300d7fe63, /* 1358 */
128'h8082450180820007802345050103b783, /* 1359 */
128'h8f999201020596130103b7830083b703, /* 1360 */
128'h059b00c6f5638e9dfff706930003b703, /* 1361 */
128'he6630103b70340a786bb87aa9d9dfff7, /* 1362 */
128'hb823001706938082852e0007002300b6, /* 1363 */
128'h4881bfe900d7002307850007c68300d3, /* 1364 */
128'h06100693488540a0053be68100055663, /* 1365 */
128'h385986ba4e250ff6f81304100693c219, /* 1366 */
128'h046e67630ff3751302b6733b0005061b, /* 1367 */
128'h8fa306850ff5751302b6563b0305051b, /* 1368 */
128'he9630300051340e685bbfe718532fea6, /* 1369 */
128'h068500f6802302d007930008876302f5, /* 1370 */
128'h86ba2581000680230015559b40e6853b, /* 1371 */
128'hbf5d00a8053b808200b61b63fff5081b, /* 1372 */
128'h178240c807bbb7d92585fea68fa30685, /* 1373 */
128'h802326050006c8830007c30397ba9381, /* 1374 */
128'h011cf0ca7119b7f10685011780230066, /* 1375 */
128'he0dafc86e4d6e8d2eccef4a6f8a2597d, /* 1376 */
128'h02500993f82af02ef42afc3e843684b2, /* 1377 */
128'h77a277420209591303000a9306c00a13, /* 1378 */
128'h178276820017079bc52d8f1d0004c503, /* 1379 */
128'h0201039304850135086304d7ff639381, /* 1380 */
128'h048905450f630014c503bfe1e7bff0ef, /* 1381 */
128'hfd07879bcb9d0004c783035510634781, /* 1382 */
128'h0014c503478100f6f36346a50ff7f793, /* 1383 */
128'h069302a6eb6306d50f63064006930489, /* 1384 */
128'hf55d08f509630630079304d50f630580, /* 1385 */
128'h6b066aa66a4669e6790674a6744670e6, /* 1386 */
128'hb74d048d0024c503808261090007051b, /* 1387 */
128'h0700071300a76c6306e50e6307300713, /* 1388 */
128'ha00d46014685003800840b13f6e51ee3, /* 1389 */
128'hf6e510e30780071302e5006307500713, /* 1390 */
128'h001636134685003800840b13fa850613, /* 1391 */
128'hb693003800840b13f8b50693a81145c1, /* 1392 */
128'h0005059be37ff0ef400845a946010016, /* 1393 */
128'h00044503a809ddbff0ef002802010393, /* 1394 */
128'hb5fd845ad93ff0ef00840b1302010393, /* 1395 */
128'h4db010ef852201247433600000840b13, /* 1396 */
128'hf436715db7f18522020103930005059b, /* 1397 */
128'hf0efe436e4c6e0c2fc3ef83aec061034, /* 1398 */
128'h862ef436f032715d8082616160e2e8df, /* 1399 */
128'he4c6e0c2fc3ef83aec06100005931014, /* 1400 */
128'hf62e710d8082616160e2e69ff0efe436, /* 1401 */
128'hee060808100005931234862afe36fa32, /* 1402 */
128'he3fff0efe436eec6eac2e6bee2baea22, /* 1403 */
128'h6135645260f28522129020ef0808842a, /* 1404 */
128'h8302000303630087b303679c691c8082, /* 1405 */
128'h47170205979304b7ee63479d80824501, /* 1406 */
128'hec061101439c97ba83f96c2707130000, /* 1407 */
128'hf55c08c52483795c878297bae426e822, /* 1408 */
128'h02f457b39381020497930c5010ef7540, /* 1409 */
128'h7d5c808261054501e91c64a2644260e2, /* 1410 */
128'h659c95aa058e05e135f1bfd9617cbfe9, /* 1411 */
128'he406e02211418082557d8082557db7e9, /* 1412 */
128'hb303679c681c00055e63ff5ff0ef842a, /* 1413 */
128'h8302014160a264028522000307630207, /* 1414 */
128'h47ad8082557d80820141640260a24501, /* 1415 */
128'h817564a7879300004797150200a7eb63, /* 1416 */
128'h80828ca505130000651780826108953e, /* 1417 */
128'h102347a1715d83020007b303679c691c, /* 1418 */
128'he83ee42e078517824785d23e47d502f1, /* 1419 */
128'hf0efcc3ed402e486100c200007930030, /* 1420 */
128'hfe63400407374d148082616160a6fd3f, /* 1421 */
128'h230134032381308345018082450100e6, /* 1422 */
128'h3823dc01011380822401011322813483, /* 1423 */
128'h3c232291342385a2980101f104132281, /* 1424 */
128'h0a04c703f579f95ff0ef1a0534832211, /* 1425 */
128'h0dd447830dd4c70302f71c630a044783, /* 1426 */
128'h02f710630c0447830c04c70302f71663, /* 1427 */
128'h0593461100f71a630e0447830e04c703, /* 1428 */
128'hfb600513d55156f010ef0d4485130d44, /* 1429 */
128'h20eff4063e800513842af0227179b761, /* 1430 */
128'hc202c40200011023858a460185226ea0, /* 1431 */
128'h6cc020ef7d000513e509842af21ff0ef, /* 1432 */
128'h10234785717980826145740270a28522, /* 1433 */
128'hc195842ac402c23ef406f022478500f1, /* 1434 */
128'h8ff9f80787934ad4008007b745386914, /* 1435 */
128'h8fd98f55400006b78f75600006b78ff5, /* 1436 */
128'h47b2e119ec9ff0ef8522858a4601c43e, /* 1437 */
128'h102347b5711d80826145740270a2c43c, /* 1438 */
128'hf852fc4ee0ca07c55783c23e47d500f1, /* 1439 */
128'he4a6e8a26a056989fdf949370107979b, /* 1440 */
128'h080909134495c43e842e8aaaec86f456, /* 1441 */
128'hf0ef8556858a4601e00a0a13e0098993, /* 1442 */
128'h0135f7b3c7891005f79345b2ed0de73f, /* 1443 */
128'h051300005517c78d0125f7b305479363, /* 1444 */
128'h64a6644660e6fba00513d4bff0ef7265, /* 1445 */
128'hc6e334fd808261257aa27a4279e26906, /* 1446 */
128'h3e80051300f057630014079b347dfe04, /* 1447 */
128'h00005517fc8049e34501b7555d8020ef, /* 1448 */
128'h2783bf7df9200513d09ff0ef6fc50513, /* 1449 */
128'h47d5c42e00f1102347c17139e7a919c5, /* 1450 */
128'hf0efc23e842af426fc06f822858a4601, /* 1451 */
128'h46014495cb918b891b842783c11dde3f, /* 1452 */
128'h70e2f8ed34fdc901dcdff0ef8522858a, /* 1453 */
128'h80824501bfd545018082612174a27442, /* 1454 */
128'h84b6892a4785e8a2ec86e0cae4a6711d, /* 1455 */
128'h260102f1102302c9270347c906d7f663, /* 1456 */
128'h0030cc3ee42e4755d432cf3108c92783, /* 1457 */
128'hd75ff0efc83eca26d23a854a100c4785, /* 1458 */
128'h02f1102347b10497f0634785e529842a, /* 1459 */
128'hd55ff0efd23ed402854a100c47f54601, /* 1460 */
128'h8522c43ff0ef6565051300005517c11d, /* 1461 */
128'hbf6147c580826125690664a6644660e6, /* 1462 */
128'hb7c54401b7d50004841bb74d02f6063b, /* 1463 */
128'he456e852ec4ef04af426f822fc067139, /* 1464 */
128'h482010ef8ab684b28a2e4148842ace05, /* 1465 */
128'h4d638cbfa0ef852200b44583c11d892a, /* 1466 */
128'h0000551700b67a63014485b368100005, /* 1467 */
128'h08c92583a0894481bd9ff0ef60c50513, /* 1468 */
128'he4030109378389a6f96decdff0ef854a, /* 1469 */
128'h854a85d6865286a2844e0089f3630207, /* 1470 */
128'h408989b308c96783fc851ae3f01ff0ef, /* 1471 */
128'h744270e2fc0999e39aa2028784339a22, /* 1472 */
128'h808261216aa26a4269e274a279028526, /* 1473 */
128'h0086969bc23e47f500f1102347997139, /* 1474 */
128'hf426f8228ed10106161b8edd030007b7, /* 1475 */
128'hf0ef8526858a4601440dc43684aafc06, /* 1476 */
128'h70e2d91ff0ef85263e800593e919c53f, /* 1477 */
128'h4d18bfcdfc79347d8082612174a27442, /* 1478 */
128'h34239fb923213823bffc07b7db010113, /* 1479 */
128'h07372331342322913c23248130232411, /* 1480 */
128'h85a2980101f104131ce7f56349013ffc, /* 1481 */
128'h1a04b7831e051863892ac09ff0ef84aa, /* 1482 */
128'hb5031aa4b023766020ef20000513e799, /* 1483 */
128'h123010ef85a2200006131e0503631a04, /* 1484 */
128'h0713000047171cf76b6347210c044783, /* 1485 */
128'h1ff78793400407b753b897ba078a1f67, /* 1486 */
128'h8007071367050d44278300e7fd63cc98, /* 1487 */
128'h0a044783f8dc00d773630147d69307a6, /* 1488 */
128'he7810019f9938b8506f48f2309b44983, /* 1489 */
128'h8a6308f480a30b344783c7890e244783, /* 1490 */
128'h8fa309c44783c7898b890a0447830009, /* 1491 */
128'h07c60c848613091407130e24478306f4, /* 1492 */
128'he0fc07c6468109d405130a844783fcdc, /* 1493 */
128'h0105959b0087979b00074583fff74783, /* 1494 */
128'h00098c634685c39197aeffe745839fad, /* 1495 */
128'h02b787b30dd4478302f585b30e044583, /* 1496 */
128'h04098f63fca714e30621070de21c07ce, /* 1497 */
128'h171b0107979b468508d4470308e44783, /* 1498 */
128'h07330e04470397ba08c447039fb90087, /* 1499 */
128'h4783f8fc07ce02e787b30dd4478302f7, /* 1500 */
128'h9fb90107171b0187979b08a4470308b4, /* 1501 */
128'h9fb9088447039fb90087171b08944703, /* 1502 */
128'h8b850a044783f4fc07a6c319f4fc54d8, /* 1503 */
128'h06134685ce81e3918bfd09c44783c789, /* 1504 */
128'h07a34785ed35e0bff0ef852645850af0, /* 1505 */
128'h979bc7b98b850e0446830af447830af4, /* 1506 */
128'h278300098663c79954dc08f4aa2300a6, /* 1507 */
128'h86bb00a6969b0dd44783f8dc07a60d44, /* 1508 */
128'h308308f480230a74478308d4ac2302f6, /* 1509 */
128'h2301390323813483854a240134032481, /* 1510 */
128'h00a7d71b50fc80822501011322813983, /* 1511 */
128'h02f707bb278527058bfd8b7d0057d79b, /* 1512 */
128'h20efd1691a04b503892abf4d08f4aa23, /* 1513 */
128'hbf455929bf555951bf651a04b0235c80, /* 1514 */
128'h229134232281382322113c23dc010113, /* 1515 */
128'h468102b7e16302f58863478923213023, /* 1516 */
128'h39038526230134032381308354a9c585, /* 1517 */
128'hffc5879b808224010113228134832201, /* 1518 */
128'h45850b900613842e4685fef760e34705, /* 1519 */
128'h99f5ffe4059bf57184aad1fff0ef892a, /* 1520 */
128'hf0ef854a85a2980101f10413f1e92581, /* 1521 */
128'hb75ddf400493f7d50b944783e51998df, /* 1522 */
128'hf022f406e44ee84aec267179b74d84aa, /* 1523 */
128'h892e9be10079f6930ff5f99308154783, /* 1524 */
128'hc519cc7ff0ef84aa45850b3006138edd, /* 1525 */
128'h852685ca00091c6300f51e63842a57b5, /* 1526 */
128'h013505a315e010ef8526842a875ff0ef, /* 1527 */
128'h8082614569a2694264e2740270a28522, /* 1528 */
128'h289134232881382328113c23d6010113, /* 1529 */
128'h275134232741382327313c2329213023, /* 1530 */
128'h259134232581382325713c2327613023, /* 1531 */
128'h4d180ac7e963478923b13c2325a13023, /* 1532 */
128'h87933ffc07b79f3dbff7879bbffc07b7, /* 1533 */
128'h210505130000551784ae8b32892abfe7, /* 1534 */
128'h5517e7b90016779307e9460300e7eb63, /* 1535 */
128'h8522f8400413f96ff0ef232505130000, /* 1536 */
128'h28013903288134832901340329813083, /* 1537 */
128'h26013b0326813a8327013a0327813983, /* 1538 */
128'h24013d0324813c8325013c0325813b83, /* 1539 */
128'h55170989270380822a01011323813d83, /* 1540 */
128'h060a81630045aa83db4520a505130000, /* 1541 */
128'hcb8902ecf7bb0005ac83e79102eaf7bb, /* 1542 */
128'hbf415429f24ff0ef2105051300005517, /* 1543 */
128'h009c9c9be3994b8502eadabb02c92783, /* 1544 */
128'h4e114e85478189d6856200c488138c0a, /* 1545 */
128'h00030d6302e8f33b0017859b00082883, /* 1546 */
128'h4c81b7c1ee4ff0ef2085051300005517, /* 1547 */
128'h80630065202302e8d33bb7f14b814a81, /* 1548 */
128'h96bbcb898b850107c78397a6078e0208, /* 1549 */
128'h0821013309bb0ffbfb9300dbebb300be, /* 1550 */
128'h55178a09000b8963fbc596e387ae0511, /* 1551 */
128'h7a1302f10a13f00600e31ea505130000, /* 1552 */
128'hee0519e3842af94ff0ef854a85d2fe0a, /* 1553 */
128'h0087979b0106161b09ea478309fa4603, /* 1554 */
128'h551785ce01367a63963e09da47839e3d, /* 1555 */
128'h0084c783b5c1e56ff0ef1da505130000, /* 1556 */
128'hf9938b89c71989b60017f7130a7a4683, /* 1557 */
128'h059b4611450547010016e993c3990fe6, /* 1558 */
128'h001878130017581b4b189726070e0017, /* 1559 */
128'h0187979b0027571b00b517bb02080463, /* 1560 */
128'hc70d4189d99b4187d79b8b050189999b, /* 1561 */
128'h8263fcc592e3872e0ff9f99300f9e9b3, /* 1562 */
128'h051300005517ef898b850a6a478302d9, /* 1563 */
128'h00f9f9b3fff7c793b591370020ef18e5, /* 1564 */
128'h051300005517cb898b8509ba4783bfd1, /* 1565 */
128'h4783e20b02e3b51d547ddbaff0ef1be5, /* 1566 */
128'h854a45850af006134685e3958b850afa, /* 1567 */
128'h0e0a47830afa07a34785e569a21ff0ef, /* 1568 */
128'h0d934d010880049308f92a2300a7979b, /* 1569 */
128'h854a458586260ff6f69301acd6bb08c0, /* 1570 */
128'h92e32d210ff4f4932485ed499f1ff0ef, /* 1571 */
128'h0ff6f693019ad6bb08f00d134c81ffb4, /* 1572 */
128'hf4932485e9359cbff0ef854a45858626, /* 1573 */
128'h8aa609b00d934d61ffa492e32ca10ff4, /* 1574 */
128'hf6930196d6bb45858656000c26834c81, /* 1575 */
128'hfa932ca12a85e13999dff0ef854a0ff6, /* 1576 */
128'h98e30c110ff4f493248dffac90e30ffa, /* 1577 */
128'h975ff0ef854a458509c0061386defdb4, /* 1578 */
128'h01379b630a7a4783d4fb0de34785ed19, /* 1579 */
128'h842a957ff0ef854a458509b006134685, /* 1580 */
128'h945ff0ef854a45850a70061386cebb3d, /* 1581 */
128'hf0ef842ae406e0221141b32ddd79842a, /* 1582 */
128'h07630187b303679c681c00055e63810f, /* 1583 */
128'h60a245058302014160a2640285220003, /* 1584 */
128'hf04af822fc06f4267139808201416402, /* 1585 */
128'h04f592635529478500f5866384aa4791, /* 1586 */
128'h4955842e07c4d78300f1102303700793, /* 1587 */
128'hf0efc43ec24a8526858a46010107979b, /* 1588 */
128'h1f634791c24a00f110234799ed19d52f, /* 1589 */
128'hd34ff0ef8526858a4601c43e478900f4, /* 1590 */
128'h14e3478580826121790274a2744270e2, /* 1591 */
128'h00f5f3634f5c6918ee09b7cdc402fef4, /* 1592 */
128'h0007059b00e7f46385be27814f1887ae, /* 1593 */
128'h691c80828082c2cff06f02c50823dd0c, /* 1594 */
128'hf4a6fc86f8a2070d4b9c711910000737, /* 1595 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 1596 */
128'h679c681cc509f11ff0ef842ac17c8fd9, /* 1597 */
128'hfd0505130000551702042423eb8d6b9c, /* 1598 */
128'h79068526744670e6f8500493bacff0ef, /* 1599 */
128'h7ca27c427be26b066aa66a4669e674a6, /* 1600 */
128'h478df93ff0eff3e54481541c80826109, /* 1601 */
128'h852202042c2302f4082347851af42c23, /* 1602 */
128'h8522681c421010ef7d000513ba2ff0ef, /* 1603 */
128'h2e2308842783f94584aa97826b9c679c, /* 1604 */
128'h8522d85c478508f422231a0428231804, /* 1605 */
128'h8522f1dff0ef852245814601b72ff0ef, /* 1606 */
128'h05a345d000ef8522f14984aacf2ff0ef, /* 1607 */
128'h4bdc00ff8737681c00f1102347a10005, /* 1608 */
128'h460147d50aa00713e3991aa007138ff9, /* 1609 */
128'h4703e911bf8ff0efc23ec43a8522858a, /* 1610 */
128'hcc1c800207b700f715630aa0079300c1, /* 1611 */
128'h4b0502900a934a55037009933e900913, /* 1612 */
128'h858a460140000cb780020c3700ff8bb7, /* 1613 */
128'he13dbb6ff0efc402c252013110238522, /* 1614 */
128'h0177f7b3c25a4bdc015110234c18681c, /* 1615 */
128'h858a4601c43e0197e7b301871563c43e, /* 1616 */
128'h397d0007ca6347b2ed1db8eff0ef8522, /* 1617 */
128'h4c14bf45331010ef3e80051306090863, /* 1618 */
128'hc43ccc188001073700e6856380020737, /* 1619 */
128'h0ca3478506041e23d45c8b8541e7d79b, /* 1620 */
128'hf0ef852202f51f63f9200793b55d18f4, /* 1621 */
128'hd663443ced09c34ff0ef85224581c04f, /* 1622 */
128'hf0ef85224585bfd118f40c2347850007, /* 1623 */
128'ha10ff0efe4c5051300005517d965c1cf, /* 1624 */
128'hf3227161551cb58584aab595fa100493, /* 1625 */
128'hf6defadafed6e352e74eeb4aef26f706, /* 1626 */
128'h45018baae3b54401e6eeeaeaeee6f2e2, /* 1627 */
128'h8ca3198bc783c7b1199bc7831ff010ef, /* 1628 */
128'h008c479d460104f110234789e7b5180b, /* 1629 */
128'h120500e3842aabaff0efc482c2be855e, /* 1630 */
128'h855e008c46014495cf818b851b8ba783, /* 1631 */
128'ha423f4fd34fd100503e3842aaa0ff0ef, /* 1632 */
128'h8522d55d842ad99ff0ef855ea031020b, /* 1633 */
128'h7b567af66a1a69ba695a64fa741a70ba, /* 1634 */
128'ha7838082615d6db66d566cf67c167bb6, /* 1635 */
128'hb16ff0ef855e0407c163180b8c23048b, /* 1636 */
128'h3e80091390810205149316d010ef4501, /* 1637 */
128'h048ba783f155842ab36ff0ef855e4585, /* 1638 */
128'h051312a96ee3149010ef85260007cc63, /* 1639 */
128'h00fbac23400007b7bfe91d7010ef0640, /* 1640 */
128'h478502fba6238b8541e7d79b048ba783, /* 1641 */
128'h1ee345111aa60f63450dbf0506fb9e23, /* 1642 */
128'h4006061b40010637a029400406370ea6, /* 1643 */
128'h8993000049978a9d0036d61b00cbac23, /* 1644 */
128'ha6830f86460396ce964e068a8a3d8069, /* 1645 */
128'h00c7d61b02d606bb018ba88345051086, /* 1646 */
128'ha42304cba823180bae231a0ba8238a05, /* 1647 */
128'h00d5183b8abd0107d69b08dba22308db, /* 1648 */
128'h02cba683090ba8231408dc63090ba623, /* 1649 */
128'h0107571b003f06b70107979b14068e63, /* 1650 */
128'h97b3070907854721938117828fd98ff5, /* 1651 */
128'hb4230c0bb0230a0bbc23030787b300e7, /* 1652 */
128'hb8230e0bb0230c0bbc230c0bb8230c0b, /* 1653 */
128'ha70308fba6230107d463200007930afb, /* 1654 */
128'hc21508fba82300e7f46320000793090b, /* 1655 */
128'h0107979b471100e78e63577d04cba783, /* 1656 */
128'hf0efc282c4be04e11023855e008c4601, /* 1657 */
128'h4601495507cbd78304f11023479d902f, /* 1658 */
128'h8e4ff0efc4bec2ca855e008c0107979b, /* 1659 */
128'h80a357fd08fbaa234785e40516e3842a, /* 1660 */
128'h855ee2051ae3842ac9aff0ef855e08fb, /* 1661 */
128'h842affbfe0ef855e00b545830f7000ef, /* 1662 */
128'h100007b754075a63018ba703e0051fe3, /* 1663 */
128'hd78306f110230370079304fba0232789, /* 1664 */
128'hd4bed2ca855e0107979b108c460107cb, /* 1665 */
128'h07930bf104934905d2caed05880ff0ef, /* 1666 */
128'h4a11d48206f11023988102091a930330, /* 1667 */
128'hd05aec56e826855e108c08104b210a85, /* 1668 */
128'hbb45842afe0a16e33a7dc131850ff0ef, /* 1669 */
128'h0165d59bbd9940030637a7a940020637, /* 1670 */
128'h16f16685b54d08bba82300b515bb89bd, /* 1671 */
128'h571b17828fd501e7569b8ff50027979b, /* 1672 */
128'h569b00ff05374098b5558b1d938100f7, /* 1673 */
128'h569b8e698fd50087161b0187179b0187, /* 1674 */
128'h27818fd58ef1f00706138fd167410087, /* 1675 */
128'h8ecd0187169b0187559b40d804fbaa23, /* 1676 */
128'h8f558f718ecd0087571b8de90087159b, /* 1677 */
128'h4689212700638b3d0187d71b04ebac23, /* 1678 */
128'h02d7971300ebac238001073720d70263, /* 1679 */
128'ha0238fd920000737040ba78300075963, /* 1680 */
128'h57971ef71863800107b7018ba70304fb, /* 1681 */
128'hf0be4d05040ba903639c232787930000, /* 1682 */
128'h6204849300003497020d1a13044ba783, /* 1683 */
128'hfe07fc1383f979130ff1079300f97933, /* 1684 */
128'h278100f977b300e797bb478540980a05, /* 1685 */
128'h109c840b0b1b4a81017d8b3716078563, /* 1686 */
128'h0197f7b300f977b340dc0007ac8397d6, /* 1687 */
128'h07b700fc8d6345a1400007b714078163, /* 1688 */
128'h40bc85b3100005b700fc886345912000, /* 1689 */
128'h0e051c638daa971ff0ef855e0015b593, /* 1690 */
128'h47912000073700ec8d6347a140000737, /* 1691 */
128'h001cb79340fc8cb3100007b700ec8863, /* 1692 */
128'h01a78663409cdfdfe0ef855e02fbaa23, /* 1693 */
128'h47d50af1102347994d850ce79163470d, /* 1694 */
128'hd53e00fde7b317c12d81810007b7d33e, /* 1695 */
128'hc93ee552e162855e110c040007930110, /* 1696 */
128'h09b794638bbd010c4783e941e91fe0ef, /* 1697 */
128'h17ed088ba58314079a631afba823409c, /* 1698 */
128'h855e460118fbae2308bba2230017b793, /* 1699 */
128'h03700793fe07fd930ff10793947ff0ef, /* 1700 */
128'h0107979b4601475507cbd7830af11023, /* 1701 */
128'he35fe0efd53ee03ad33a8cee855e110c, /* 1702 */
128'h4791d502d33a0af1102347b56702e915, /* 1703 */
128'he552e16ee43e855e110c011004000713, /* 1704 */
128'h670267a20e050c63e0dfe0efe03ac93a, /* 1705 */
128'ha2231afba823017d85b74785f3ed37fd, /* 1706 */
128'hf0ef855e840585934601180bae23096b, /* 1707 */
128'h0000379704a1eafa94e347a10a918c9f, /* 1708 */
128'h9285051300005517e6f49fe349c78793, /* 1709 */
128'h071b80011737b61ddf400413cbdfe0ef, /* 1710 */
128'h0307971300ebac2380020737b519a007, /* 1711 */
128'h0ff104934905bbc580030737de075ee3, /* 1712 */
128'h3a7d09053ac54a159881190201000ab7, /* 1713 */
128'h1030c33e47d508f110234799020a0863, /* 1714 */
128'hdc3ef84af426c556855e010c04000793, /* 1715 */
128'hfbe18b8583a54cdcd0051ce3d61fe0ef, /* 1716 */
128'h0087d79b0087961bf006869366c144dc, /* 1717 */
128'hda06d9e3040ba70302e796938fd18ff5, /* 1718 */
128'h68e34581472db35d04fba02300876793, /* 1719 */
128'hb54511872583974e837902079713eaf7, /* 1720 */
128'ha783f006869300ff0537040d859366c1, /* 1721 */
128'h961b8f510187971b0187d61b0d91000d, /* 1722 */
128'hae238fd98ff58f510087d79b8e690087, /* 1723 */
128'h00c7579b46a5008ca703fdb59ee3fefd, /* 1724 */
128'h1c63800306b7018ba60300f6f8638bbd, /* 1725 */
128'ha78397b6078a2ee686930000369704d6, /* 1726 */
128'h67c100cca68308fbae230087171b1487, /* 1727 */
128'h27810126d71b8fd10186d61b8ff917fd, /* 1728 */
128'h02e6073b3e800613c305c38d03f77713, /* 1729 */
128'ha02302d606bb02f757bb8a8d0106d69b, /* 1730 */
128'ha7831afbaa231b0ba7830adba2230afb, /* 1731 */
128'h08fba82308fba62320000793c79919cb, /* 1732 */
128'ha7030005062300051523484000ef855e, /* 1733 */
128'h8693aaa78793ccccd6b7aaaab7b708cb, /* 1734 */
128'h37b3068600d036b327818ef98ff9ccc6, /* 1735 */
128'h36b38ef90f068693f0f0f6b79fb500f0, /* 1736 */
128'h8ef9f0068693ff0106b79fb5068a00d0, /* 1737 */
128'h8f750207161376c19fb5068e00d036b3, /* 1738 */
128'h92010a8bb783d11c9fb9071200e03733, /* 1739 */
128'hc603074bd68307abd70302c7d7b3ed10, /* 1740 */
128'h02450513764585930000459784aa06fb, /* 1741 */
128'h077bc883070ba803a95fe0effef53623, /* 1742 */
128'h0188569b0108571b0088579b06cbc603, /* 1743 */
128'h459726810ff777130ff878130ff7f793, /* 1744 */
128'ha603a5ffe0ef04d48513742585930000, /* 1745 */
128'h569b0624851373e5859300004597074b, /* 1746 */
128'h8526a3ffe0ef8a3d8abd0146561b0106, /* 1747 */
128'h100007b7b8d102fba42347857e4010ef, /* 1748 */
128'h6ce31a0bb683400407b704fba0232785, /* 1749 */
128'h0737bb956bc5051300004517e691ecf7, /* 1750 */
128'hf6930c46c78304fba0230017079b7000, /* 1751 */
128'h00c7f693ce910027f6931adba42303f7, /* 1752 */
128'h6713040ba70304eba0230217071bc689, /* 1753 */
128'he793040ba783c7998b8504eba0230107, /* 1754 */
128'ha583044ba783040baa0304fba02300c7, /* 1755 */
128'h84930000349700fa7a33855e4601088b, /* 1756 */
128'h1b0b0b1300003b174a85db4ff0ef19e4, /* 1757 */
128'h00fa97bb409c1e2c8c9300003c974c2d, /* 1758 */
128'h1909091300003917cbb5278100fa77b3, /* 1759 */
128'h17ed00494703409c10000db720000d37, /* 1760 */
128'h77b30009270340dc04f718630017b793, /* 1761 */
128'h45850b70061300894683c3a18ff900fa, /* 1762 */
128'h06134681c131debfe0ef855e0fb6f693, /* 1763 */
128'ha823088ba783ddbfe0ef855e45850b70, /* 1764 */
128'h855e035baa2308fba223180bae231a0b, /* 1765 */
128'hf7649fe304a1fb9911e30931973fe0ef, /* 1766 */
128'h2783bb6d925fe0ef5905051300004517, /* 1767 */
128'h8663471100d789634721400006b70009, /* 1768 */
128'h855e02ebaa230017b71341b787b301a7, /* 1769 */
128'h2683f941808ff0ef855e408c933fe0ef, /* 1770 */
128'hef8d1afba823409ce79d0046f7930089, /* 1771 */
128'hae2308bba2230017b79317ed088ba583, /* 1772 */
128'h9fdfe0ef855ecb0ff0ef855e460118fb, /* 1773 */
128'h855e45850b7006130ff6f693bb91fd31, /* 1774 */
128'h9713fcfc65e34581b7c9f521d31fe0ef, /* 1775 */
128'h00ec4641bf6d11872583974e83790207, /* 1776 */
128'hd78304f11023478d6da000ef06cb8513, /* 1777 */
128'h47d5855ec4be0107979b008c460107cb, /* 1778 */
128'h018ba783ec051b63842a96ffe0efc2be, /* 1779 */
128'h102347a506fb9e2304e157830007d663, /* 1780 */
128'h979b008c460107cbd783c2be479d04f1, /* 1781 */
128'hea051163842a93bfe0efc4be855e0107, /* 1782 */
128'h04dbae23018ba50345e6475647c646b6, /* 1783 */
128'h4000063706bba42306eba22306fba023, /* 1784 */
128'h8ca602e345098a3d01a6d61bf2c51a63, /* 1785 */
128'h061b40010637f0a609634505f0c54363, /* 1786 */
128'hc56ce54ff06ffa100413f0eff06f2006, /* 1787 */
128'h18b50d238082557d8082557d80824501, /* 1788 */
128'h1141ef9d439cde278793000057978082, /* 1789 */
128'hdcf7262300005717842ae406e0224785, /* 1790 */
128'h852200055563aeefe0ef852212a000ef, /* 1791 */
128'h0dc000ef13e000ef02c00513fc5ff0ef, /* 1792 */
128'h571780824501808201414501640260a2, /* 1793 */
128'h114102e790636394631cd9a707130000, /* 1794 */
128'hf60fe0efe40653e505130000451785aa, /* 1795 */
128'h04630fc7a60380820141853e478160a2, /* 1796 */
128'hec06110141488082853ebfd187b600a6, /* 1797 */
128'h006365a210354703c105fbdff0efe42e, /* 1798 */
128'h60e200f70c630ff007930815470302b7, /* 1799 */
128'h45018082610560e25535eb3fe06f6105, /* 1800 */
128'he822ec06e4261101bfcdf8400513bfe5, /* 1801 */
128'he501cf0ff0ef842acd09f7dff0ef84ae, /* 1802 */
128'h8082610564a2644260e2e0800f840413, /* 1803 */
128'h071b4388b847879300005797bfd55535, /* 1804 */
128'h0000579780820f8505138082c3980015, /* 1805 */
128'h879300005797110180824388b6c78793, /* 1806 */
128'h0094176384beec06e4266380e822cce7, /* 1807 */
128'hc78119a447838082610564a2644260e2, /* 1808 */
128'h879300005797b7d56000a9cff0ef8522, /* 1809 */
128'h8082b207a12300005797e79ce39cc9e7, /* 1810 */
128'he11ce7886798c867879300005797e508, /* 1811 */
128'h849300005497e4a6711d8082e308e518, /* 1812 */
128'hec5ef05af456f852fc4e6080e8a2c6e4, /* 1813 */
128'h00004a1789aae0caec86e06ae466e862, /* 1814 */
128'h00004b1741ca8a9300004a9742ca0a13, /* 1815 */
128'h00050c1b424b8b9300004b97424b0b13, /* 1816 */
128'h6446029415634d29a08c8c9300004c97, /* 1817 */
128'h6be27b027aa27a4279e2690664a660e6, /* 1818 */
128'h612557250513000045176d026ca26c42, /* 1819 */
128'hc36389524c1cc7914901541cddcfe06f, /* 1820 */
128'he0ef638c855a0fc42603681c89560007, /* 1821 */
128'h601cdb2fe0ef855e85ca00090663dbef, /* 1822 */
128'h01a98863da4fe0ef856685e200978e63, /* 1823 */
128'hb771600032a010ef9905051300004517, /* 1824 */
128'h4d1cc1414401e04ae426ec06e8221101, /* 1825 */
128'hc7bd651ccbad511ccbbd4d5ccfad4401, /* 1826 */
128'h10ef45051c00059384aa892ec7ad639c, /* 1827 */
128'h0ef52c234799c57c57fdcd21842a2000, /* 1828 */
128'h0405282303253023e90410f502a34785, /* 1829 */
128'h16f43c2391c78793fffff797e65ff0ef, /* 1830 */
128'h0000179718f430232be7879300001797, /* 1831 */
128'h85220ea42e23681c18f434232ae78793, /* 1832 */
128'h60e28522e99ff0ef10f400230247c783, /* 1833 */
128'h56971bc0106f80826105690264a26442, /* 1834 */
128'h02d786b365186294611c8aa686930000, /* 1835 */
128'h836d8f3d0127d713e118973600176713, /* 1836 */
128'h8d5d00f717bb40f007b300f7553b93ed, /* 1837 */
128'hfc3ff06fae4505130000551780822501, /* 1838 */
128'hfe9ff0ef842afefff0efe022e4061141, /* 1839 */
128'h808201412501640260a28d410105151b, /* 1840 */
128'h14020005041bfdbff0efe022e4061141, /* 1841 */
128'h0141640260a28d4115029001fd1ff0ef, /* 1842 */
128'hfee78fa30785fff5c703058587aa8082, /* 1843 */
128'hc703058500c7896387aa962a8082fb75, /* 1844 */
128'hc70387aa8082fb65fee78fa30785fff5, /* 1845 */
128'h0785fff5c7030585eb09001786930007, /* 1846 */
128'he21987aab7d587b68082fb75fee78fa3, /* 1847 */
128'h963efb7d001786930007c70387b68082, /* 1848 */
128'he291fed70fa300178713fff5c6830585, /* 1849 */
128'hb7cd87ba8082000780a300c715638082, /* 1850 */
128'h979b40f707bbfff5c783000547030585, /* 1851 */
128'h8082853ef37d0505e3994187d79b0187, /* 1852 */
128'h000547030585a839478100c59463962e, /* 1853 */
128'h4187d79b0187979b40f707bbfff5c783, /* 1854 */
128'h47830ff5f5938082853eff790505e399, /* 1855 */
128'h4501bfcd0505c399808200b793630005, /* 1856 */
128'h808200b79363000547830ff5f5938082, /* 1857 */
128'h8533e7010007c70387aabfcd0505dffd, /* 1858 */
128'h842ae42ee8221101bfcd0785808240a7, /* 1859 */
128'h47830ff5f593952265a2fe5ff0efec06, /* 1860 */
128'h60e24501fe857be3157d00b786630005, /* 1861 */
128'hc70300b7856387aa95aa808261056442, /* 1862 */
128'h862ab7fd0785808240a78533e7010007, /* 1863 */
128'h0fe38082ea9940c785330007c68387aa, /* 1864 */
128'hb7d50785fe081be3000748030705fed8, /* 1865 */
128'h40d785330007c60387aa86aabfcd872e, /* 1866 */
128'h1be300074803070500c80a638082ea11, /* 1867 */
128'h00054703bff90785bfd5872e8082fe08, /* 1868 */
128'h0007c6830785fee68fe380824501eb19, /* 1869 */
128'he426e8221101bfd587aeb7e50505fafd, /* 1870 */
128'h8e07879300005797e519842a84aeec06, /* 1871 */
128'h4783942af9dff0ef85a68522cc116380, /* 1872 */
128'h852244018c07b22300005797ef810004, /* 1873 */
128'hf0ef852285a68082610564a2644260e2, /* 1874 */
128'h050500050023c78100054783c519f9ff, /* 1875 */
128'h6104e4261101bfd988a7bc2300005797, /* 1876 */
128'hc501f73ff0ef8526842ac891e822ec06, /* 1877 */
128'h64a28526644260e2e008050500050023, /* 1878 */
128'hc68387aacf9900054783c11d80826105, /* 1879 */
128'h00e780238082e3110017c703ce810007, /* 1880 */
128'h0075779380824501b7e5078900d780a3, /* 1881 */
128'h8fd507a2808204c79063963e87aacb9d, /* 1882 */
128'h40e88833469d00c508b3872aff6d377d, /* 1883 */
128'h078e02e787335761003657930106ef63, /* 1884 */
128'h0721bfd10ff5f6934725bfc1963a97aa, /* 1885 */
128'h0a63bf6dfeb78fa30785bfe1fef73c23, /* 1886 */
128'h9e63963e87aacb9d8b9d00a5e7b300b5, /* 1887 */
128'hff07bc2307a1ff8738030721808202c7, /* 1888 */
128'h07b357e100365713ff06e8e340f88833, /* 1889 */
128'h872ebfc100e507b3963e95ba070e02f7, /* 1890 */
128'hfff5c7030585bfe1469d00c508b387aa, /* 1891 */
128'h852e842af0227179bf65fee78fa30785, /* 1892 */
128'h6622dcdff0efe02ee84af406e432ec26, /* 1893 */
128'hfff6091300c564636582892ace1184aa, /* 1894 */
128'h70a200040023f79ff0ef944a864a8522, /* 1895 */
128'he02211418082614564e2694285267402, /* 1896 */
128'h60a28522f57ff0ef00a5e963842ae406, /* 1897 */
128'h40b6073300c506b395b2808201416402, /* 1898 */
128'h802316fd0005c78315fdd7e500e587b3, /* 1899 */
128'h8082853e478100c51563962ab7fd00f6, /* 1900 */
128'h05850505fbed9f990005c70300054783, /* 1901 */
128'h8de300054783808200c51363962ab7dd, /* 1902 */
128'hec26852e842af0227179bfc50505feb7, /* 1903 */
128'h0005049bd1fff0ef89aee84af406e44e, /* 1904 */
128'h00995b630005091bd13ff0ef8522c889, /* 1905 */
128'h614569a2694264e2740270a285224401, /* 1906 */
128'hd175f8bff0ef397d852285ce86268082, /* 1907 */
128'h450100c514630ff5f593962abfe90405, /* 1908 */
128'h853efeb70be300150793000547038082, /* 1909 */
128'h87aa260100c7ef630ff5f59347c1b7ed, /* 1910 */
128'hfeb71ce30007c7038082853e4781e601, /* 1911 */
128'h873b47a1c31d00757713b7f5367d0785, /* 1912 */
128'hfcb81ce30007c80387aa0007069b40e7, /* 1913 */
128'h8e1d953e938102071793faf5078536fd, /* 1914 */
128'h96938fd90107179300b7e73300859793, /* 1915 */
128'h8a1deb1187aa27018edd003657130207, /* 1916 */
128'hbfcd367d0785f8b71fe30007c703d24d, /* 1917 */
128'h0007c70300d80a63008785130007b803, /* 1918 */
128'h377d87aabfa5fef51be30785f8b712e3, /* 1919 */
128'h11630300079300054703e7a9419cb7f1, /* 1920 */
128'h86b32ea78793000027970015470308f7, /* 1921 */
128'h77130207071bc6898a850006c68300e7, /* 1922 */
128'h97ba0025470304d71b63078006930ff7, /* 1923 */
128'h4198c19c47c1c3b10447f7930007c783, /* 1924 */
128'h1663030007930005470302f71c6347c1, /* 1925 */
128'h973e29a70713000027170015478302f7, /* 1926 */
128'h0ff7f7930207879bc7098b0500074703, /* 1927 */
128'hbf7d47a18082050900e7936307800713, /* 1928 */
128'hc632ec06006c842ee8221101bf6d47a9, /* 1929 */
128'h081300002817468100c16583f63ff0ef, /* 1930 */
128'h460300f806330007079b000547032568, /* 1931 */
128'h644260e2ec0500089863044678930006, /* 1932 */
128'h879b00088b6300467893808261058536, /* 1933 */
128'hb7d196be050502d586b3feb7f4e3fd07, /* 1934 */
128'hfc97879b0ff7f793fe07079bc6098a09, /* 1935 */
128'hf04afc06f426f8227139b7e1e008b7cd, /* 1936 */
128'h65a2b0dff0ef84b2842ae42e00063023, /* 1937 */
128'h80826121790274a2744270e25529e901, /* 1938 */
128'h82e367e2f5dff0ef8522082c892a862e, /* 1939 */
128'hfd279be307858f81cb010007c703fe87, /* 1940 */
128'h00054683b7e94501e088fcf718e347a9, /* 1941 */
128'h05051141f2dff06f00e6846302d00713, /* 1942 */
128'h8082014140a0053360a2f23ff0efe406, /* 1943 */
128'h0693601cf0dff0ef842ee406e0221141, /* 1944 */
128'h069300e6ea6302d704630007c70304b0, /* 1945 */
128'h069380820141640260a202d70e630470, /* 1946 */
128'hc683fed716e306b0069302d7076304d0, /* 1947 */
128'h0027c683fce69fe3052a069007130017, /* 1948 */
128'h052ab7e9e01c078d00e6986304200713, /* 1949 */
128'h006c842ee8221101bfd50789bff1052a, /* 1950 */
128'h2817468100c16583e0fff0efc632ec06, /* 1951 */
128'h06330007079b00054703102808130000, /* 1952 */
128'hec0500089863044678930006460300f8, /* 1953 */
128'h8b6300467893808261058536644260e2, /* 1954 */
128'h050502d586b3feb7f4e3fd07879b0008, /* 1955 */
128'h0ff7f793fe07079bc6098a09b7d196be, /* 1956 */
128'he406e0221141b7e1e008b7cdfc97879b, /* 1957 */
128'h0007c70304b00693601cf87ff0ef842e, /* 1958 */
128'h02d70e630470069300e6ea6302d70463, /* 1959 */
128'h02d7076304d0069380820141640260a2, /* 1960 */
128'h069007130017c683fed716e306b00693, /* 1961 */
128'h9863042007130027c683fce69fe3052a, /* 1962 */
128'h0789bff1052a052ab7e9e01c078d00e6, /* 1963 */
128'h95bff0efe589842ae406e0221141bfd5, /* 1964 */
128'h0287879300002797fff5c70300a405b3, /* 1965 */
128'h60a2e7198b1100074703973efff58513, /* 1966 */
128'h4703fea47ae3157d80820141557d6402, /* 1967 */
128'h60a26402f77d8b1100074703973e0005, /* 1968 */
128'hf06f4581d7dff06f0141050545814629, /* 1969 */
128'h550300a10723812100a107a31141fa5f, /* 1970 */
128'h639c4ba78793000047978082014100e1, /* 1971 */
128'h4781aa5ff06f95be9201160291811582, /* 1972 */
128'h069b8082853ee3190005470345a94625, /* 1973 */
128'h9fb902f587bb00d667630ff6f693fd07, /* 1974 */
128'h842ee406e0221141bff90505fd07879b, /* 1975 */
128'h02b455bb45a900b7f86347a500a04563, /* 1976 */
128'h60a2640202a4753b4529fe7ff0ef357d, /* 1977 */
128'h07e2081007935000006f030505130141, /* 1978 */
128'h44f730230000471744f7302300004717, /* 1979 */
128'he4264324041300004417e82211018082, /* 1980 */
128'h600ca15ff0efec06600885aa84ae862e, /* 1981 */
128'h11018082610564a26442e00c95a660e2, /* 1982 */
128'h849300004497e4264087879300004797, /* 1983 */
128'h9b050513000045176380e82260903f64, /* 1984 */
128'hc0ef85a26088b87fd0ef85a29c11ec06, /* 1985 */
128'h9a85051300004517862286aa608ce63f, /* 1986 */
128'hb61fd0ef9b45051300004517b6dfd0ef, /* 1987 */
128'h00055e6384ff90efef65051300000517, /* 1988 */
128'h05130000451740a005b364a260e26442, /* 1989 */
128'h610564a260e26442b39fd06f61059a65, /* 1990 */
128'h870fa0ef8432e406e02211416680006f, /* 1991 */
128'h450180820141640260a2557d00850363, /* 1992 */
128'h852289aae64e01258413f22271698082, /* 1993 */
128'h04b30505f7eff0ef892eea4aee26f606, /* 1994 */
128'he93ff0ef95260505f72ff0ef852600a4, /* 1995 */
128'h0000479704e7ee631ff00793fff5071b, /* 1996 */
128'h0000351784aaf50ff0ef852230a7ae23, /* 1997 */
128'hf2630ff007939526f42ff0ef71c50513, /* 1998 */
128'h051300003517842af32ff0ef852204a7, /* 1999 */
128'h05130000451700a405b3f24ff0ef6fe5, /* 2000 */
128'h69b2695264f2741270b2a8bfd0ef9165, /* 2001 */
128'h2cf72023000047172000079380826155, /* 2002 */
128'h3597863ff0ef850a458110000613b755, /* 2003 */
128'h01294703deaff0ef850a6ba585930000, /* 2004 */
128'h8e8585930000459700f7096302f00793, /* 2005 */
128'h4797df2ff0ef850a85a2dfaff0ef850a, /* 2006 */
128'h051300004517858a439027a787930000, /* 2007 */
128'h4717451107e208100793a1bfd0ef8ce5, /* 2008 */
128'hf0ef26f731230000471726f731230000, /* 2009 */
128'hd77ff0ef450102a79f2300004797d85f, /* 2010 */
128'h859300004597461102a7992300004797, /* 2011 */
128'h1123000047174785eb1ff0ef854e0265, /* 2012 */
128'h478de04ae426ec06e8221101b79122f7, /* 2013 */
128'hd37ff0ef84ae450d892a08c7df638432, /* 2014 */
128'h55030000451708a7956325010004d783, /* 2015 */
128'h06a79a6325010024d783d21ff0ef1f25, /* 2016 */
128'hf0ef4511dabff0ef00448513ffc4059b, /* 2017 */
128'h550300004517faa79f2300004797d05f, /* 2018 */
128'hfaa79523000047974611cf1ff0ef1c25, /* 2019 */
128'h4535e2bff0ef854afa05859300004597, /* 2020 */
128'hf0ef45151985d58300004597256000ef, /* 2021 */
128'h879300004797240000ef02000513d1bf, /* 2022 */
128'h16f71a230000471727850007d7831827, /* 2023 */
128'h0087cf63278d439c1687879300004797, /* 2024 */
128'h60e26442905fd0ef7d85051300003517, /* 2025 */
128'h64a2644260e2d49ff06f6105690264a2, /* 2026 */
128'h0105c783f022f4067179808261056902, /* 2027 */
128'h578300f10f230115c78300f10fa34709, /* 2028 */
128'h70a2740202e78a63470d00e78e6301e1, /* 2029 */
128'h842a8b3fd06f61457b85051300003517, /* 2030 */
128'h85228a3fd0efe42e7905051300003517, /* 2031 */
128'h41907402d8bff06f614570a265a27402, /* 2032 */
128'h3823dc010113ebfff06f614505c170a2, /* 2033 */
128'h893284ae842a23213023229134232281, /* 2034 */
128'he60ff0ef22113c230028218006134581, /* 2035 */
128'hea2ff0efe802c44a08282040061385a6, /* 2036 */
128'h2301340323813083f63ff0ef8522002c, /* 2037 */
128'h47978082240101132201390322813483, /* 2038 */
128'h8593000045974611cb8107e7d7830000, /* 2039 */
128'h504000efe40611418082cf3ff06fe665, /* 2040 */
128'h27051001a70300e57763878e1041e703, /* 2041 */
128'h150260a21007e78310a7a22310e1a023, /* 2042 */
128'h110180824501808201418d5d91011782, /* 2043 */
128'h00ef842afc1ff0ef84aae426e822ec06, /* 2044 */
128'h60e29101150202f407b33e8007934400, /* 2045 */
128'h11418082610564a28d0502a7d5336442, /* 2046 */
128'h47b7414000ef842af95ff0efe022e406, /* 2047 */
128'h1502640260a202f407b324078793000f, /* 2048 */
128'he822ec061101808202a7d53301419101, /* 2049 */
128'h3e2000ef892af63ff0ef84aae04ae426, /* 2050 */
128'h0285543324040413000f443702a48533, /* 2051 */
128'h644260e2fe856ee3f45ff0ef0405944a, /* 2052 */
128'h009894b7e426110180826105690264a2, /* 2053 */
128'hf363892268048493842ae04aec06e822, /* 2054 */
128'hf47dfa1ff0ef41240433854a89260084, /* 2055 */
128'h00b5002380826105690264a2644260e2, /* 2056 */
128'h0147c503410007b78082000545038082, /* 2057 */
128'hf7930147478341000737808202057513, /* 2058 */
128'h8223410007b7808200a70023dfe50207, /* 2059 */
128'h00e78023476d00e78623f80007130007, /* 2060 */
128'h8423fc70071300e78623470d00078223, /* 2061 */
128'he0221141808200e788230200071300e7, /* 2062 */
128'h0141640260a2e50900044503842ae406, /* 2063 */
128'h879300002797b7f50405fa5ff0ef8082, /* 2064 */
128'h0007470397aa973e811100f57713f4e7, /* 2065 */
128'h1101808200f5802300e580a30007c783, /* 2066 */
128'h4503fd1ff0efec068121842a002ce822, /* 2067 */
128'h002cf5dff0ef00914503f65ff0ef0081, /* 2068 */
128'hf4bff0ef00814503fb7ff0ef0ff47513, /* 2069 */
128'h80826105644260e2f43ff0ef00914503, /* 2070 */
128'h54e14461892af406e84aec26f0227179, /* 2071 */
128'h4503f81ff0ef0ff57513002c0089553b, /* 2072 */
128'hf0bff0ef00914503f13ff0ef34610081, /* 2073 */
128'h80826145694264e2740270a2fe9410e3, /* 2074 */
128'h03800413892af406e84aec26f0227179, /* 2075 */
128'hf3fff0ef0ff57513002c0089553354e1, /* 2076 */
128'hf0ef00914503ed1ff0ef346100814503, /* 2077 */
128'h6145694264e2740270a2fe9410e3ec9f, /* 2078 */
128'h00814503f13ff0efec06002c11018082, /* 2079 */
128'h610560e2e9fff0ef00914503ea7ff0ef, /* 2080 */
128'hf8227139439c02678793000047978082, /* 2081 */
128'h856384b2842e892aec4efc06f04af426, /* 2082 */
128'h2501f3afb0efdce505130000451702b7, /* 2083 */
128'h74a2744270e2fea7ad2300004797c10d, /* 2084 */
128'h2f230000471757fd8082612169e27902, /* 2085 */
128'hd98505130000451785ca86260074fcf7, /* 2086 */
128'hfca7a22300004797c50d2501814fb0ef, /* 2087 */
128'h430505130000351785a6049675634632, /* 2088 */
128'hb775faf72323000047174785d0cfd0ef, /* 2089 */
128'h37970009099b00c4591be05ff0ef4521, /* 2090 */
128'h00094503993e0039791342a787930000, /* 2091 */
128'h47979c25bf5d320010ef854ede7ff0ef, /* 2092 */
128'h842a85aae0221141bf95f687a5230000, /* 2093 */
128'h100fcb2fd0efe4064005051300003517, /* 2094 */
128'h60a264028322f14025730ff0000f0000, /* 2095 */
128'h4605114183020141db05859300002597, /* 2096 */
128'hf2850513000045170e85859300003597, /* 2097 */
128'h00003517c9112501d79fa0efe022e406, /* 2098 */
128'h3517c62fd06f014160a264023e450513, /* 2099 */
128'h000035974605c56fd0ef3f2505130000, /* 2100 */
128'hd9bfa0efcac505130000451740458593, /* 2101 */
128'h3517b7e13fc5051300003517c5112501, /* 2102 */
128'h051300000517c26fd0ef27a505130000, /* 2103 */
128'ha72300004797ea07ad2300004797e985, /* 2104 */
128'h0000479700054863842a904f90efea07, /* 2105 */
128'h60a26402408005b3cf81439cea078793, /* 2106 */
128'h4517be2fd06f01412505051300003517, /* 2107 */
128'h3517c5112501b9afb0efc42505130000, /* 2108 */
128'h8593000035974605bfb93aa505130000, /* 2109 */
128'h00003517c5112501cb9fa0ef450101e5, /* 2110 */
128'h00000023ee1ff0ef8522b7813a450513, /* 2111 */
128'h4537a001d69ff0efe406250111419002, /* 2112 */
128'h0000471780824501808224050513000f, /* 2113 */
128'h0017869300756513157d631ce1470713, /* 2114 */
128'h06338082953e055e10d00513e3089536, /* 2115 */
128'hfd1ff0efe4328532ec06e822110102b5, /* 2116 */
128'h60e28522944ff0ef45816622c509842a, /* 2117 */
128'h05130000351711418082808261056442, /* 2118 */
128'hee5fc0ef42000537b28fd0efe40633e5, /* 2119 */
128'h808245018082450180820141450160a2, /* 2120 */
128'h87361141808202f5553347a9b0002573, /* 2121 */
128'he40632a505130000351785aa862e86b2, /* 2122 */
128'he0221141a001cbbff0ef4505aecfd0ef, /* 2123 */
128'h9522408007b3f57ff0efe406952e842a, /* 2124 */
128'h450580824505808201418d7d640260a2, /* 2125 */
128'h842ef406ec26f0227179808245058082, /* 2126 */
128'h450164e2740270a20096186300c684bb, /* 2127 */
128'h6622e37fc0efe432852285b280826145, /* 2128 */
128'h8082450980824509bff9260520040413, /* 2129 */
128'h45018082450180828082808280824509, /* 2130 */
128'h4781e426e822ec061101bbbff06f8082, /* 2131 */
128'h00c7986300d5043300d584b300379693, /* 2132 */
128'h0004380380826105450164a2644260e2, /* 2133 */
128'h0513000035176090600c02e803636098, /* 2134 */
128'h05130000351785a28626a2afd0ef29e5, /* 2135 */
128'he0ca711dbf5d0785a001a1afd0ef2b65, /* 2136 */
128'hf852fc4ee8a22b65051300003517892a, /* 2137 */
128'h8b2ee466e4a6ec86e862ec5ef05af456, /* 2138 */
128'h3b972a2a0a1300003a179eafd0ef4401, /* 2139 */
128'h0c1300003c17fff949932aab8b930000, /* 2140 */
128'h85e600040c9b9c6fd0ef85524ac12aec, /* 2141 */
128'h855203649863448187ca9bafd0ef855e, /* 2142 */
128'h458187ca9a4fd0ef856285e69acfd0ef, /* 2143 */
128'h051300003517fd5417e3040502b49b63, /* 2144 */
128'h8a85008486b3a889450198afd0ef2d65, /* 2145 */
128'h6398e39840e9873300349713c689873e, /* 2146 */
128'h873e8a856390008586b3bf5d07a10485, /* 2147 */
128'h058e02e60d6340e9873300359713c689, /* 2148 */
128'h00003517944fd0ef2385051300003517, /* 2149 */
128'h64a6644660e6557d938fd0ef26450513, /* 2150 */
128'h6ca26c426be27b027aa27a4279e26906, /* 2151 */
128'hfc56e0d27159bfa507a1058580826125, /* 2152 */
128'hf45ef85ae4ceeca6020005138aaa6a05, /* 2153 */
128'h8b2ee46ee86aec66e8caf0a2f486f062, /* 2154 */
128'h3c179c4a0a134981b3fff0ef44818bb2, /* 2155 */
128'h0cb300fa8db30034979359ac0c130000, /* 2156 */
128'hd0ef232505130000351703749b6300fb, /* 2157 */
128'h7c027ba26a0669a6694670a674068bef, /* 2158 */
128'h85567b4264e685da86266da26d426ce2, /* 2159 */
128'he0ef842abddfe0efe33ff06f61657ae2, /* 2160 */
128'hf7b3bcbfe0ef892abd1fe0ef8d2abd7f, /* 2161 */
128'h643300a96533010d1d1b0105151b0344, /* 2162 */
128'hb02300acb0238d4191011402150201a4, /* 2163 */
128'h0039f7930985aadff0ef4521ef8100ad, /* 2164 */
128'h7139b7ad0485a9dff0ef0007c50397e2, /* 2165 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2166 */
128'hb69fe0ef892ab6ffe0ef842ab75fe0ef, /* 2167 */
128'h8d450109179b0105151bb63fe0ef84aa, /* 2168 */
128'h47818d5d9101178265a2660215028fc1, /* 2169 */
128'h744200c79c63974e00e5883300379713, /* 2170 */
128'hf06f6121863e69e2854e790274a270e2, /* 2171 */
128'h8f2900083703e3148ea907856314d79f, /* 2172 */
128'hf822fc06e032e42e7139b7f100e83023, /* 2173 */
128'he0ef842aafdfe0ef89aaec4ef04af426, /* 2174 */
128'h151baebfe0ef84aaaf1fe0ef892aaf7f, /* 2175 */
128'h65a2660215028fc18d450109179b0105, /* 2176 */
128'h00e588330037971347818d5d91011782, /* 2177 */
128'h854e790274a270e2744200c79c63974e, /* 2178 */
128'h8e8907856314d01ff06f6121863e69e2, /* 2179 */
128'h7139b7f100e830238f0900083703e314, /* 2180 */
128'h89aaec4ef04af426f822fc06e032e42e, /* 2181 */
128'ha79fe0ef892aa7ffe0ef842aa85fe0ef, /* 2182 */
128'h8d450109179b0105151ba73fe0ef84aa, /* 2183 */
128'h47818d5d9101178265a2660215028fc1, /* 2184 */
128'h744200c79c63974e00e5883300379713, /* 2185 */
128'hf06f6121863e69e2854e790274a270e2, /* 2186 */
128'h00083703e31402a686b307856314c89f, /* 2187 */
128'he032e42e7139b7e100e8302302a70733, /* 2188 */
128'ha09fe0ef89aaec4ef04af426f822fc06, /* 2189 */
128'he0ef84aa9fdfe0ef892aa03fe0ef842a, /* 2190 */
128'h15028fc18d450109179b0105151b9f7f, /* 2191 */
128'h0037971347818d5d9101178265a26602, /* 2192 */
128'h74a270e2744200c79c63974e00e58833, /* 2193 */
128'he111c0dff06f6121863e69e2854e7902, /* 2194 */
128'h00083703e31402a6d6b3078563144505, /* 2195 */
128'he032e42e7139b7d100e8302302a75733, /* 2196 */
128'h989fe0ef89aaec4ef04af426f822fc06, /* 2197 */
128'he0ef84aa97dfe0ef892a983fe0ef842a, /* 2198 */
128'h15028fc18d450109179b0105151b977f, /* 2199 */
128'h0037971347818d5d9101178265a26602, /* 2200 */
128'h74a270e2744200c79c63974e00e58833, /* 2201 */
128'h6314b8dff06f6121863e69e2854e7902, /* 2202 */
128'h00e830238f4900083703e3148ec90785, /* 2203 */
128'hf04af426f822fc06e032e42e7139b7f1, /* 2204 */
128'h892a90bfe0ef842a911fe0ef89aaec4e, /* 2205 */
128'h179b0105151b8fffe0ef84aa905fe0ef, /* 2206 */
128'h9101178265a2660215028fc18d450109, /* 2207 */
128'h9c63974e00e588330037971347818d5d, /* 2208 */
128'h863e69e2854e790274a270e2744200c7, /* 2209 */
128'h3703e3148ee907856314b15ff06f6121, /* 2210 */
128'he032e42e7139b7f100e830238f690008, /* 2211 */
128'h899fe0ef89aaec4ef04af426f822fc06, /* 2212 */
128'he0ef84aa88dfe0ef892a893fe0ef842a, /* 2213 */
128'h14828fc18cc90109179b0105151b887f, /* 2214 */
128'h0037169347018fc59081178265a26602, /* 2215 */
128'h74a270e2744200c71c6396ae00d98833, /* 2216 */
128'h0533a9dff06f6121863a69e2854e7902, /* 2217 */
128'he8ca7159bfc9070500a83023e28800f7, /* 2218 */
128'he0d2e4cef0a2d965051300003517892a, /* 2219 */
128'h89aeec66eca6f486f062f45ef85afc56, /* 2220 */
128'hd80a0a1300003a17cc9fc0ef44018b32, /* 2221 */
128'hd90c0c1300003c17d88b8b9300003b97, /* 2222 */
128'h85a2fff44493ca7fc0ef855204000a93, /* 2223 */
128'h14fd460140900cb3c99fc0ef8885855e, /* 2224 */
128'h85520566186397ce00f905b300361793, /* 2225 */
128'h6622c73fc0ef856285a2c7bfc0efe432, /* 2226 */
128'h1be32405e12984aaa03ff0ef854a85ce, /* 2227 */
128'h70a6c53fc0efd9e5051300003517fb54, /* 2228 */
128'h7b427ae26a0669a664e6694685267406, /* 2229 */
128'h876600167693808261656ce27c027ba2, /* 2230 */
128'hbfc154fdbf590605e198e3988726c291, /* 2231 */
128'hf0a2cc2505130000351784aaeca67159, /* 2232 */
128'hec66f062f45ef85afc56e0d2e4cee8ca, /* 2233 */
128'h3997bf3fc0ef44018ab2892ee86af486, /* 2234 */
128'h3b97faab0b1300003b17caa989930000, /* 2235 */
128'h3c97ca2c0c1300003c17faab8b930000, /* 2236 */
128'hbc1fc0ef854e04000a13caac8c930000, /* 2237 */
128'hc0ef856285a2000bbd03cba500147793, /* 2238 */
128'h00f485b300361793fffd45134601baff, /* 2239 */
128'h85a2b93fc0efe432854e05561c6397ca, /* 2240 */
128'h91bff0ef852685ca6622b8bfc0ef8566, /* 2241 */
128'h051300003517fb441ae32405e5298d2a, /* 2242 */
128'h694664e6856a740670a6b6bfc0efcb65, /* 2243 */
128'h6d426ce27c027ba27b427ae26a0669a6, /* 2244 */
128'h876a00167693bf49000b3d0380826165, /* 2245 */
128'hb7e15d7db7790605e198e398872ac291, /* 2246 */
128'he4a6bd25051300003517842ae8a2711d, /* 2247 */
128'hfc4eec86e862ec5ef05af456f852e0ca, /* 2248 */
128'h091300003917b07fc0ef4c018ab284ae, /* 2249 */
128'h8b9300003b97bc6b0b1300003b17bbe9, /* 2250 */
128'h000c099bae5fc0ef854a10000a13bceb, /* 2251 */
128'h010c1793008c1713ad9fc0ef855a85ce, /* 2252 */
128'h020c17138fd9018c17130187e7b38fd9, /* 2253 */
128'h17138fd9030c17138fd9028c17138fd9, /* 2254 */
128'h972600e406b30036171346018fd9038c, /* 2255 */
128'h855e85cea95fc0efe432854a05561763, /* 2256 */
128'h89aa81dff0ef852285a66622a8dfc0ef, /* 2257 */
128'hbb85051300003517f94c19e30c05e91d, /* 2258 */
128'h79e2690664a6854e644660e6a6dfc0ef, /* 2259 */
128'he31c808261256c426be27b027aa27a42, /* 2260 */
128'h84aaf4a67119bff159fdb74d0605e29c, /* 2261 */
128'he8d2eccef0caf8a2ae85051300003517, /* 2262 */
128'hec6efc86f06af466f862fc5ee0dae4d6, /* 2263 */
128'h0a1300003a17a17fc0ef44018b32892e, /* 2264 */
128'h498507f00b93ad6c8c9300003c97acea, /* 2265 */
128'h08000a93ad4d0d1300003d1703f00c13, /* 2266 */
128'h873b9e3fc0ef856685a29ebfc0ef8552, /* 2267 */
128'h003617934601008995b300e99733408b, /* 2268 */
128'hc0efe432855205661a6397ca00f486b3, /* 2269 */
128'h852685ca66229b7fc0ef856a85a29bff, /* 2270 */
128'h3517fb541be32405e1398daaf46ff0ef, /* 2271 */
128'h856e744670e6997fc0efae2505130000, /* 2272 */
128'h7c427be26b066aa66a4669e6790674a6, /* 2273 */
128'he38c008c6663808261096de27d027ca2, /* 2274 */
128'hb7f15dfdbfe5e298e398bf610605e28c, /* 2275 */
128'hf8a2a02505130000351784aaf4a67119, /* 2276 */
128'hf466f862fc5ee0dae4d6e8d2eccef0ca, /* 2277 */
128'h931fc0ef44018b32892eec6efc86f06a, /* 2278 */
128'h9f0c8c9300003c979e8a0a1300003a17, /* 2279 */
128'h0d1300003d1703f00c13498507f00b93, /* 2280 */
128'h856685a2905fc0ef855208000a939eed, /* 2281 */
128'h008996b300f997b3408b87bb8fdfc0ef, /* 2282 */
128'h85b3003617134601fff6c693fff7c793, /* 2283 */
128'h8d1fc0efe432855205661a63974a00e4, /* 2284 */
128'hf0ef852685ca66228c9fc0ef856a85a2, /* 2285 */
128'h00003517fb5417e32405e1398daae58f, /* 2286 */
128'h74a6856e744670e68a9fc0ef9f450513, /* 2287 */
128'h7ca27c427be26b066aa66a4669e67906, /* 2288 */
128'he194e314008c6663808261096de27d02, /* 2289 */
128'h7119b7f15dfdbfe5e19ce31cbf610605, /* 2290 */
128'hf0caf8a2914505130000351784aaf4a6, /* 2291 */
128'hf06af466f862fc5ee0dae4d6e8d2ecce, /* 2292 */
128'h3997843fc0ef44018a32892eec6efc86, /* 2293 */
128'h0a93902c0c1300003c178fa989930000, /* 2294 */
128'h00003c9703f00b9308100b134d0507f0, /* 2295 */
128'hc0ef856285a2817fc0ef854e8fcc8c93, /* 2296 */
128'h173300fd17b3408b07bb408a873b80ff, /* 2297 */
128'h008d16b300fd17b30024079b8f5d00ed, /* 2298 */
128'h003616934601fff7c313fff748938fd5, /* 2299 */
128'hc0efe432854e05461c6396ca00d48533, /* 2300 */
128'h852685ca6622fc6fc0ef856685a2fcef, /* 2301 */
128'h1be3080007932405ed298daad56ff0ef, /* 2302 */
128'h70e6fa2fc0ef8ee5051300003517f8f4, /* 2303 */
128'h6b066aa66a4669e6790674a6856e7446, /* 2304 */
128'h7813808261096de27d027ca27c427be2, /* 2305 */
128'he28c85be00081363859a008bea630016, /* 2306 */
128'hbfc585bafe081be385c6b7610605e10c, /* 2307 */
128'h051300002517892af0ca7119bf755dfd, /* 2308 */
128'hfc86ec6ef06af466fc5ee8d2ecce7fe5, /* 2309 */
128'h4b81e03289aef862e0dae4d6f4a6f8a2, /* 2310 */
128'h00002c977e4a0a1300002a17f2cfc0ef, /* 2311 */
128'h47854da17f4d0d1300002d177ecc8c93, /* 2312 */
128'hf00fc0ef85524401003b949b01779c33, /* 2313 */
128'hfffc4a93ef4fc0ef856685da00848b3b, /* 2314 */
128'h1063974e00e908330036171367824601, /* 2315 */
128'hc0ef856a85daed6fc0efe432855206f6, /* 2316 */
128'he9318b2ac5eff0ef854a85ce6622ecef, /* 2317 */
128'h90e3040007932b85fbb41be38c562405, /* 2318 */
128'h70e6ea2fc0ef7ee5051300002517fafb, /* 2319 */
128'h6b066aa66a4669e6790674a6855a7446, /* 2320 */
128'h7513808261096de27d027ca27c427be2, /* 2321 */
128'h060500b83023e30c85d6e11185e20016, /* 2322 */
128'h84aaf4cef8cafca67175b7e95b7db749, /* 2323 */
128'he4dee8daecd6f0d2698502000513892e, /* 2324 */
128'h4a81e032f46ef86ae122e506fc66e0e2, /* 2325 */
128'h899332ac0c1300003c174a01892ff0ef, /* 2326 */
128'h4d818bca8b26ae6c8c9300003c979c49, /* 2327 */
128'h866e04fd956396da003d969367824d21, /* 2328 */
128'h020a0863ed45842aba2ff0ef852685ca, /* 2329 */
128'h60aa8522df4fc0ef7685051300002517, /* 2330 */
128'h6ba66b466ae67a0679a6794674e6640a, /* 2331 */
128'h8b4a4a05808261497da27d427ce26c06, /* 2332 */
128'h908fe0ef842a90efe0efec36b7758ba6, /* 2333 */
128'h664267a28fcfe0efe42a902fe0efe82a, /* 2334 */
128'h140215028c510106161b8d5d0105151b, /* 2335 */
128'he28828a7b523000037978d4166e29101, /* 2336 */
128'h078500fb86330006c683018786b34781, /* 2337 */
128'h033df7b3ffa795e300d600230ff6f693, /* 2338 */
128'h8a9b001a879bfbdfe0ef4521ef910ba1, /* 2339 */
128'h0d85fa9fe0ef0007c50397e68b8d0007, /* 2340 */
128'h892af0d2f4cef8ca7175bfa1547dbf0d, /* 2341 */
128'he4dee8daecd6fca66a050200051389ae, /* 2342 */
128'h4b018cb2f46ee122e506f86afc66e0e2, /* 2343 */
128'h0a1321248493000034974a81f73fe0ef, /* 2344 */
128'h4d818c4e8bca9c6d0d1300003d179c4a, /* 2345 */
128'h866e059d956397de00fc06b3003d9793, /* 2346 */
128'h020a8863e579842aa82ff0ef854a85ce, /* 2347 */
128'h60aa8522cd4fc0ef6485051300002517, /* 2348 */
128'h6ba66b466ae67a0679a6794674e6640a, /* 2349 */
128'h8bce4a85808261497da27d427ce26c06, /* 2350 */
128'hd0ef842afedfd0efe836ec3eb7758c4a, /* 2351 */
128'h6622fdbfd0efe02afe1fd0efe42afe7f, /* 2352 */
128'h15028c518d590106161b0105151b6702, /* 2353 */
128'h67e216a7b923000037978d4191011402, /* 2354 */
128'h00f6902393c117c20004d783e38866c2, /* 2355 */
128'h0044d78300f6912393c117c20024d783, /* 2356 */
128'h93c117c20064d78300f6922393c117c2, /* 2357 */
128'he87fe0ef4521ef91034df7b300f69323, /* 2358 */
128'h0007c50397ea8b8d00078b1b001b079b, /* 2359 */
128'h80826505b789547dbf290d85e73fe0ef, /* 2360 */
128'h842afca6e122fff586138932f8ca7175, /* 2361 */
128'hf4ce56a505130000251785aa962a84ae, /* 2362 */
128'hf46ef86afc66e0e2e4dee8daecd6f0d2, /* 2363 */
128'h0014d9930044d793bd8fc0efec36e506, /* 2364 */
128'h2b1744854a81e43e99a20034d793e83e, /* 2365 */
128'h2c17552b8b9300002b97552b0b130000, /* 2366 */
128'h2d17552c8c9300002c97552c0c130000, /* 2367 */
128'h3a1755ad8d9300002d9755ad0d130000, /* 2368 */
128'h0513000025170299786306aa0a130000, /* 2369 */
128'h794674e68556640a60aab7afc0ef54e5, /* 2370 */
128'h7d427ce26c066ba66b466ae67a0679a6, /* 2371 */
128'h0663b52fc0ef855a85a6808261497da2, /* 2372 */
128'hb40fc0ef8562b46fc0ef855e85ca0009, /* 2373 */
128'h920ff0ef852265a2b38fc0ef856a85e6, /* 2374 */
128'h49636762010a2783b28fc0ef856eed15, /* 2375 */
128'h4d05051300002517c58d000a358302f7, /* 2376 */
128'h9782852285ce6642008a3783b0cfc0ef, /* 2377 */
128'hb7e94a89af4fc0ef4c05051300002517, /* 2378 */
128'hbfa10485ae4fc0ef2785051300002517, /* 2379 */
128'hec26f022f4064ae50513000025177179, /* 2380 */
128'h0000251704000593c19fe0efe44ee84a, /* 2381 */
128'h4c85051300002517ab8fc0ef4ac50513, /* 2382 */
128'haa0fc0ef4ec5051300002517aacfc0ef, /* 2383 */
128'h4441a92fc0ef44852285051300002517, /* 2384 */
128'h853346054685008495b3497901f49993, /* 2385 */
128'h740270a2ff2417e3e6dff0ef24050135, /* 2386 */
128'h131b460580828082614569a2694264e2, /* 2387 */
128'h87f245a901f61e1346814881470100c5, /* 2388 */
128'h97aa0007802397aa0007802340000813, /* 2389 */
128'h13e397aa387d0007802397aa00078023, /* 2390 */
128'h26f38e15c020267302b71d632705fe08, /* 2391 */
128'h059302a68733411686b33e800513c000, /* 2392 */
128'h473302a767b302b345bb02c747334000, /* 2393 */
128'h10e39f2fc06f486505130000251702a7, /* 2394 */
128'he4061141bf51c00028f3c02026f3fac7, /* 2395 */
128'hf0ef4509f75ff0ef4505f7bff0ef4501, /* 2396 */
128'h4541f63ff0ef4521f69ff0ef4511f6ff, /* 2397 */
128'he388440007b791011502bff1f5dff0ef, /* 2398 */
128'h440007b7808225016388440007b78082, /* 2399 */
128'h7b88440007b7808225016b880007b823, /* 2400 */
128'h07b70106161b8d5d0085979b80822501, /* 2401 */
128'hef634400073747812581f7888d514400, /* 2402 */
128'hc3198b097a98440006b73e80079300b7, /* 2403 */
128'h0006e60380827388440007b7ffe537fd, /* 2404 */
128'h4785e406e0221141bfe1f71006912785, /* 2405 */
128'hf0ef250135fd0045551b00b7d863842a, /* 2406 */
128'h4503943e3fc7879300002797883dfebf, /* 2407 */
128'h07b7711da1ffe06f014160a264020004, /* 2408 */
128'h571b3006869300a7893b6685e0ca0040, /* 2409 */
128'he4a6e8a20587e7938f550089179b0189, /* 2410 */
128'hc63ec43a454d842a4589460184ae0034, /* 2411 */
128'h46010034f4dff0eff456f852fc4eec86, /* 2412 */
128'h458946010034f3fff0ef454d8a2a4589, /* 2413 */
128'h0793083886a60810f31ff0ef454d89aa, /* 2414 */
128'h00f9d8330106002300fa583355e10380, /* 2415 */
128'h060537e10107002300f5583301068023, /* 2416 */
128'hf3dff0ef854a45a1feb790e307050685, /* 2417 */
128'h1a974981874fc0ef4705051300001517, /* 2418 */
128'h10181782013407bb4a21462a8a930000, /* 2419 */
128'hf0dff0ef29854589ff07c50397ba9381, /* 2420 */
128'h051300002517ff4991e384afc0ef8556, /* 2421 */
128'h1517eefff0ef854a45a183afc0effce5, /* 2422 */
128'h00001a974981826fc0ef422505130000, /* 2423 */
128'h97a693811782013407bb4a21414a8a93, /* 2424 */
128'hb0ef8556ec1ff0ef298545890007c503, /* 2425 */
128'hb0eff825051300002517ff4992e3ffff, /* 2426 */
128'h051300001517ea3ff0ef45a1854afeff, /* 2427 */
128'h3c898993000019974481fdbfb0ef3d65, /* 2428 */
128'hc50397ba938110181782009407bb4921, /* 2429 */
128'hfb1fb0ef854ee73ff0ef24854589ff87, /* 2430 */
128'hfa1fb0eff345051300002517ff2491e3, /* 2431 */
128'h61257aa27a4279e2690664a6644660e6, /* 2432 */
128'hec56f052f44ef84afc26e0a2715d8082, /* 2433 */
128'h0a1b440184aa89328aae89aae486e85a, /* 2434 */
128'h002c054463630154053b44000b37ff86, /* 2435 */
128'h8526002c920116024089063be4dff0ef, /* 2436 */
128'h4ac133aa0a1300001a174401d9ffd0ef, /* 2437 */
128'h640660a603246863ec8b0b1300002b17, /* 2438 */
128'h808261616b426ae27a0279a2794274e2, /* 2439 */
128'h9381178200c4579b2421e0bff0ef85a6, /* 2440 */
128'hdbdff0ef852245a1b74500fb302304a1, /* 2441 */
128'h93811782009407bb4481efbfb0ef8552, /* 2442 */
128'h8552d9fff0ef248545890007c50397ce, /* 2443 */
128'h2441ed3fb0ef855aff5492e3eddfb0ef, /* 2444 */
128'hb0efe406d1450513000025171141bf61, /* 2445 */
128'h5c63badf70eff305051300000517ebff, /* 2446 */
128'hd08505130000251740a005b360a20005, /* 2447 */
128'h25179cffe06f014160a2e9bfb06f0141, /* 2448 */
128'hf822fc067139fd6fe06f21a505130000, /* 2449 */
128'hf8efe0efe05ae456e852ec4ef04af426, /* 2450 */
128'h09b74401fb4fe0ef1585051300002517, /* 2451 */
128'h013407b3449515690913000029170880, /* 2452 */
128'he41fb0ef0405854a0004059b6390078e, /* 2453 */
128'h0b1300002b174901c18f80effe9416e3, /* 2454 */
128'h2a17132a8a9300002a97440004b72f6b, /* 2455 */
128'h0007c783016907b34991142a0a130000, /* 2456 */
128'h8622240125816080608ce09c09058556, /* 2457 */
128'hb0ef25818552688c0004b823dfdfb0ef, /* 2458 */
128'h47190054579b0ff47413fd391be3deff, /* 2459 */
128'h97ba078a6cc707130000071702f76463, /* 2460 */
128'hb0ef1025051300002517878297ba439c, /* 2461 */
128'h051300002517a001929fe0ef8522dbff, /* 2462 */
128'h2517b7f5edbff0ef8522dabfb0ef0fe5, /* 2463 */
128'hbfe9ab7ff0efd97fb0ef0fa505130000, /* 2464 */
128'hc94f80efd85fb0ef0f85051300002517, /* 2465 */
128'hf0efd73fb0ef0f65051300002517b7e1, /* 2466 */
128'h000000000000000000000000bf5db8ff, /* 2467 */
128'h00000000000000000000000000000000, /* 2468 */
128'h00000000000000000000000000000000, /* 2469 */
128'h00000000000000000000000000000000, /* 2470 */
128'h00000000000000000000000000000000, /* 2471 */
128'h00000000000000000000000000000000, /* 2472 */
128'h00000000000000000000000000000000, /* 2473 */
128'h00000000000000000000000000000000, /* 2474 */
128'h00000000000000000000000000000000, /* 2475 */
128'h00000000000000000000000000000000, /* 2476 */
128'h00000000000000000000000000000000, /* 2477 */
128'h00000000000000000000000000000000, /* 2478 */
128'h00000000000000000000000000000000, /* 2479 */
128'h08082828282828080808080808080808, /* 2480 */
128'h08080808080808080808080808080808, /* 2481 */
128'h101010101010101010101010101010a0, /* 2482 */
128'h10101010101004040404040404040404, /* 2483 */
128'h01010101010101010141414141414110, /* 2484 */
128'h10101010100101010101010101010101, /* 2485 */
128'h02020202020202020242424242424210, /* 2486 */
128'h08101010100202020202020202020202, /* 2487 */
128'h00000000000000000000000000000000, /* 2488 */
128'h00000000000000000000000000000000, /* 2489 */
128'h101010101010101010101010101010a0, /* 2490 */
128'h10101010101010101010101010101010, /* 2491 */
128'h01010101010101010101010101010101, /* 2492 */
128'h02010101010101011001010101010101, /* 2493 */
128'h02020202020202020202020202020202, /* 2494 */
128'h02020202020202021002020202020202, /* 2495 */
128'hc1bdceee242070dbe8c7b756d76aa478, /* 2496 */
128'hfd469501a83046134787c62af57c0faf, /* 2497 */
128'h895cd7beffff5bb18b44f7af698098d8, /* 2498 */
128'h49b40821a679438efd9871936b901122, /* 2499 */
128'he9b6c7aa265e5a51c040b340f61e2562, /* 2500 */
128'he7d3fbc8d8a1e68102441453d62f105d, /* 2501 */
128'h455a14edf4d50d87c33707d621e1cde6, /* 2502 */
128'h8d2a4c8a676f02d9fcefa3f8a9e3e905, /* 2503 */
128'hfde5380c6d9d61228771f681fffa3942, /* 2504 */
128'hbebfbc70f6bb4b604bdecfa9a4beea44, /* 2505 */
128'h04881d05d4ef3085eaa127fa289b7ec6, /* 2506 */
128'hc4ac56651fa27cf8e6db99e5d9d4d039, /* 2507 */
128'hfc93a039ab9423a7432aff97f4292244, /* 2508 */
128'h85845dd1ffeff47d8f0ccc92655b59c3, /* 2509 */
128'h4e0811a1a3014314fe2ce6e06fa87e4f, /* 2510 */
128'heb86d3912ad7d2bbbd3af235f7537e82, /* 2511 */
128'h0c07020d08030e09040f0a05000b0601, /* 2512 */
128'h020f0c090603000d0a0704010e0b0805, /* 2513 */
128'h09020b040d060f08010a030c050e0700, /* 2514 */
128'h6c5f7465735f64735f63736972776f6c, /* 2515 */
128'h6e67696c615f64730000000000006465, /* 2516 */
128'h645f6b6c635f64730000000000000000, /* 2517 */
128'h69747465735f64730000000000007669, /* 2518 */
128'h735f646d635f6473000000000000676e, /* 2519 */
128'h74657365725f64730000000074726174, /* 2520 */
128'h6e636b6c625f64730000000000000000, /* 2521 */
128'h69736b6c625f64730000000000000074, /* 2522 */
128'h6f656d69745f6473000000000000657a, /* 2523 */
128'h655f7172695f64730000000000007475, /* 2524 */
128'h5f63736972776f6c000000000000006e, /* 2525 */
128'h00000000646d635f74726174735f6473, /* 2526 */
128'h746e695f746961775f63736972776f6c, /* 2527 */
128'h000000000067616c665f747075727265, /* 2528 */
128'h00007172695f64735f63736972776f6c, /* 2529 */
128'h695f646d635f64735f63736972776f6c, /* 2530 */
128'h5f63736972776f6c0000000000007172, /* 2531 */
128'h007172695f646e655f617461645f6473, /* 2532 */
128'h0000000087fe9e880000000087feb150, /* 2533 */
128'h004c4b40004c4b400030000020000000, /* 2534 */
128'h6d6d5f6472616f62000000020000ffff, /* 2535 */
128'h0000000087fe4ea00064637465675f63, /* 2536 */
128'h0000000087fe4d0c0000000087fe4aae, /* 2537 */
128'h00000000000000000000000000000000, /* 2538 */
128'hffffb982ffffb97effffb97effffb958, /* 2539 */
128'hffffb986ffffb986ffffb986ffffb986, /* 2540 */
128'h0000000087feb4780000000087feb468, /* 2541 */
128'h0000000087feb4a00000000087feb488, /* 2542 */
128'h0000000087feb4d00000000087feb4b8, /* 2543 */
128'h0000000087feb5000000000087feb4e8, /* 2544 */
128'h0000000087feb5300000000087feb518, /* 2545 */
128'h0000000087feb5600000000087feb548, /* 2546 */
128'h40040300400402004004010040040000, /* 2547 */
128'h40050000400405004004040140040400, /* 2548 */
128'h30000000000000030000000040050100, /* 2549 */
128'h60000000000000053000000000000001, /* 2550 */
128'h70000000000000027000000000000004, /* 2551 */
128'h00000001400000007000000000000000, /* 2552 */
128'h00000005000000012000000000000006, /* 2553 */
128'h20000000000000020000000040000000, /* 2554 */
128'h00000000100000000000000100000000, /* 2555 */
128'h1e19140f0d0c0a000000000000000000, /* 2556 */
128'h000186a00000271050463c37322d2823, /* 2557 */
128'h017d7840017d784000989680000f4240, /* 2558 */
128'h031975000319750002faf080018cba80, /* 2559 */
128'h02faf08005f5e10002faf080017d7840, /* 2560 */
128'h00000020000000000bebc2000c65d400, /* 2561 */
128'h00000200000001000000008000000040, /* 2562 */
128'h00002000000010000000080000000400, /* 2563 */
128'h0000c000000080000000600000004000, /* 2564 */
128'h37363534333231300002000000010000, /* 2565 */
128'h2043534952776f4c4645444342413938, /* 2566 */
128'h746f6f622d7520646573696d696e696d, /* 2567 */
128'h00000000647261432d445320726f6620, /* 2568 */
128'hfffff958fffff96efffff95afffff946, /* 2569 */
128'h00000000fffff992fffff958fffff980, /* 2570 */
128'he00600003800000039080000edfe0dd0, /* 2571 */
128'h00000000100000001100000028000000, /* 2572 */
128'h0000000000000000a806000059010000, /* 2573 */
128'h00000000010000000000000000000000, /* 2574 */
128'h02000000000000000400000003000000, /* 2575 */
128'h020000000f0000000400000003000000, /* 2576 */
128'h2c6874651b0000001400000003000000, /* 2577 */
128'h007665642d657261622d656e61697261, /* 2578 */
128'h2c687465260000001000000003000000, /* 2579 */
128'h0100000000657261622d656e61697261, /* 2580 */
128'h1a0000000300000000006e65736f6863, /* 2581 */
128'h313440747261752f636f732f2c000000, /* 2582 */
128'h0000003030323531313a303030303030, /* 2583 */
128'h00000000737570630100000002000000, /* 2584 */
128'h01000000000000000400000003000000, /* 2585 */
128'h000000000f0000000400000003000000, /* 2586 */
128'h40787d01380000000400000003000000, /* 2587 */
128'h03000000000000304075706301000000, /* 2588 */
128'h0300000080f0fa024b00000004000000, /* 2589 */
128'h03000000007570635b00000004000000, /* 2590 */
128'h03000000000000006700000004000000, /* 2591 */
128'h0000000079616b6f6b00000005000000, /* 2592 */
128'h7a6874651b0000001300000003000000, /* 2593 */
128'h0000766373697200656e61697261202c, /* 2594 */
128'h34367672720000000b00000003000000, /* 2595 */
128'h0b000000030000000000636466616d69, /* 2596 */
128'h0000393376732c76637369727c000000, /* 2597 */
128'h01000000850000000000000003000000, /* 2598 */
128'h6f72746e6f632d747075727265746e69, /* 2599 */
128'h04000000030000000000000072656c6c, /* 2600 */
128'h0000000003000000010000008f000000, /* 2601 */
128'h1b0000000f00000003000000a0000000, /* 2602 */
128'h000063746e692d7570632c7663736972, /* 2603 */
128'h01000000b50000000400000003000000, /* 2604 */
128'h01000000bb0000000400000003000000, /* 2605 */
128'h01000000020000000200000002000000, /* 2606 */
128'h0030303030303030384079726f6d656d, /* 2607 */
128'h6f6d656d5b0000000700000003000000, /* 2608 */
128'h67000000100000000300000000007972, /* 2609 */
128'h00000008000000000000008000000000, /* 2610 */
128'h0300000000636f730100000002000000, /* 2611 */
128'h03000000020000000000000004000000, /* 2612 */
128'h03000000020000000f00000004000000, /* 2613 */
128'h616972612c6874651b0000001f000000, /* 2614 */
128'h706d697300636f732d657261622d656e, /* 2615 */
128'h000000000300000000007375622d656c, /* 2616 */
128'h303240746e696c6301000000c3000000, /* 2617 */
128'h0d000000030000000000003030303030, /* 2618 */
128'h30746e696c632c76637369721b000000, /* 2619 */
128'hca000000100000000300000000000000, /* 2620 */
128'h07000000010000000300000001000000, /* 2621 */
128'h00000000670000001000000003000000, /* 2622 */
128'h0300000000000c000000000000000002, /* 2623 */
128'h006c6f72746e6f63de00000008000000, /* 2624 */
128'h7075727265746e690100000002000000, /* 2625 */
128'h3030634072656c6c6f72746e6f632d74, /* 2626 */
128'h04000000030000000000000030303030, /* 2627 */
128'h04000000030000000000000000000000, /* 2628 */
128'h0c00000003000000010000008f000000, /* 2629 */
128'h003063696c702c76637369721b000000, /* 2630 */
128'h03000000a00000000000000003000000, /* 2631 */
128'h0b00000001000000ca00000010000000, /* 2632 */
128'h10000000030000000900000001000000, /* 2633 */
128'h000000000000000c0000000067000000, /* 2634 */
128'he8000000040000000300000000000004, /* 2635 */
128'hfb000000040000000300000007000000, /* 2636 */
128'hb5000000040000000300000003000000, /* 2637 */
128'hbb000000040000000300000002000000, /* 2638 */
128'h75626564010000000200000002000000, /* 2639 */
128'h0000304072656c6c6f72746e6f632d67, /* 2640 */
128'h637369721b0000001000000003000000, /* 2641 */
128'h03000000003331302d67756265642c76, /* 2642 */
128'hffff000001000000ca00000008000000, /* 2643 */
128'h00000000670000001000000003000000, /* 2644 */
128'h03000000001000000000000000000000, /* 2645 */
128'h006c6f72746e6f63de00000008000000, /* 2646 */
128'h30313440747261750100000002000000, /* 2647 */
128'h08000000030000000000003030303030, /* 2648 */
128'h03000000003035373631736e1b000000, /* 2649 */
128'h00000041000000006700000010000000, /* 2650 */
128'h04000000030000000010000000000000, /* 2651 */
128'h040000000300000080f0fa024b000000, /* 2652 */
128'h040000000300000000c2010006010000, /* 2653 */
128'h04000000030000000200000014010000, /* 2654 */
128'h04000000030000000100000025010000, /* 2655 */
128'h04000000030000000200000030010000, /* 2656 */
128'h0100000002000000040000003a010000, /* 2657 */
128'h3030323440636d6d2d63736972776f6c, /* 2658 */
128'h10000000030000000000000030303030, /* 2659 */
128'h00000000000000420000000067000000, /* 2660 */
128'h14010000040000000300000000000100, /* 2661 */
128'h25010000040000000300000002000000, /* 2662 */
128'h1b0000000c0000000300000002000000, /* 2663 */
128'h0200000000636d6d2d63736972776f6c, /* 2664 */
128'h406874652d63736972776f6c01000000, /* 2665 */
128'h03000000000000003030303030303334, /* 2666 */
128'h2d63736972776f6c1b0000000c000000, /* 2667 */
128'h5b000000080000000300000000687465, /* 2668 */
128'h0400000003000000006b726f7774656e, /* 2669 */
128'h04000000030000000200000014010000, /* 2670 */
128'h06000000030000000300000025010000, /* 2671 */
128'h0300000000007fe3023e180047010000, /* 2672 */
128'h00000043000000006700000010000000, /* 2673 */
128'h01000000020000000080000000000000, /* 2674 */
128'h343440646e7277682d63736972776f6c, /* 2675 */
128'h0e000000030000000000303030303030, /* 2676 */
128'h6e7277682d63736972776f6c1b000000, /* 2677 */
128'h67000000100000000300000000000064, /* 2678 */
128'h00100000000000000000004400000000, /* 2679 */
128'h09000000020000000200000002000000, /* 2680 */
128'h2300736c6c65632d7373657264646123, /* 2681 */
128'h61706d6f6300736c6c65632d657a6973, /* 2682 */
128'h6f647473006c65646f6d00656c626974, /* 2683 */
128'h65736162656d697400687461702d7475, /* 2684 */
128'h6b636f6c630079636e6575716572662d, /* 2685 */
128'h63697665640079636e6575716572662d, /* 2686 */
128'h75746174730067657200657079745f65, /* 2687 */
128'h2d756d6d006173692c76637369720073, /* 2688 */
128'h230074696c70732d626c740065707974, /* 2689 */
128'h00736c6c65632d747075727265746e69, /* 2690 */
128'h6f72746e6f632d747075727265746e69, /* 2691 */
128'h646e6168702c78756e696c0072656c6c, /* 2692 */
128'h727265746e69007365676e617200656c, /* 2693 */
128'h6572006465646e657478652d73747075, /* 2694 */
128'h616d2c76637369720073656d616e2d67, /* 2695 */
128'h766373697200797469726f6972702d78, /* 2696 */
128'h70732d746e6572727563007665646e2c, /* 2697 */
128'h61702d747075727265746e6900646565, /* 2698 */
128'h0073747075727265746e6900746e6572, /* 2699 */
128'h6f692d6765720074666968732d676572, /* 2700 */
128'h63616d2d6c61636f6c0068746469772d, /* 2701 */
128'h0000000000000000737365726464612d, /* 2702 */
128'h0000000000203a642520656369766544, /* 2703 */
128'h00203a6425206563697665642073250a, /* 2704 */
128'h00000000203a6425206563697665440a, /* 2705 */
128'h000a656369766564206e776f6e6b6e75, /* 2706 */
128'h00000a2973252c73252870756b6f6f6c, /* 2707 */
128'h7265206c616e7265746e692070636864, /* 2708 */
128'h00000000000000000a7025202c726f72, /* 2709 */
128'h5145525f5043484420676e69646e6553, /* 2710 */
128'h4b434120504348440000000a54534555, /* 2711 */
128'h696c432050434844000000000000000a, /* 2712 */
128'h203a7373657264644120504920746e65, /* 2713 */
128'h0000000a64252e64252e64252e642520, /* 2714 */
128'h73657264644120504920726576726553, /* 2715 */
128'h0a64252e64252e64252e642520203a73, /* 2716 */
128'h6120726574756f520000000000000000, /* 2717 */
128'h252e64252e642520203a737365726464, /* 2718 */
128'h6b73616d2074654e0000000a64252e64, /* 2719 */
128'h64252e642520203a7373657264646120, /* 2720 */
128'h697420657361654c000a64252e64252e, /* 2721 */
128'h7364253a6d64253a686425203d20656d, /* 2722 */
128'h3d206e69616d6f44000000000000000a, /* 2723 */
128'h4820746e65696c4300000a2273252220, /* 2724 */
128'h000a22732522203d20656d616e74736f, /* 2725 */
128'h000000000a44455050494b53204b4341, /* 2726 */
128'h000000000000000a4b414e2050434844, /* 2727 */
128'h73657264646120646574736575716552, /* 2728 */
128'h0000000000000a646573756665722073, /* 2729 */
128'h000000000000000a732520726f727245, /* 2730 */
128'h6e6f6974706f2064656c646e61686e75, /* 2731 */
128'h656c646e61686e55000000000a642520, /* 2732 */
128'h64252065646f63706f20504348442064, /* 2733 */
128'h20676e69646e6553000000000000000a, /* 2734 */
128'h000a595245564f435349445f50434844, /* 2735 */
128'h00000000000a29732528726f72726570, /* 2736 */
128'h3a2043414d2073250000000030687465, /* 2737 */
128'h3a583230253a583230253a5832302520, /* 2738 */
128'h000a583230253a583230253a58323025, /* 2739 */
128'h484420646e65732074276e646c756f43, /* 2740 */
128'h206e6f20595245564f43534944205043, /* 2741 */
128'h00000a7325203a732520656369766564, /* 2742 */
128'h5043484420726f6620676e6974696157, /* 2743 */
128'h2020202020202020000a524546464f5f, /* 2744 */
128'h00000000000063250000000000000020, /* 2745 */
128'h0000005832302520000000000000002e, /* 2746 */
128'h00000000732573250000000000000a0a, /* 2747 */
128'h00000000007325203a646c697542202c, /* 2748 */
128'h73257a4820756c250000000000007325, /* 2749 */
128'h0000000000756c250000000000000000, /* 2750 */
128'h0073257a4863252000000000646c252e, /* 2751 */
128'h00000000007325736574794220756c25, /* 2752 */
128'h00003a786c3830250073254269632520, /* 2753 */
128'h000a73252020202000786c6c2a302520, /* 2754 */
128'h000000203a5d64255b6e6f6974636553, /* 2755 */
128'h727265207974696e6173207264646170, /* 2756 */
128'h2c7825286e666c6500000a702520726f, /* 2757 */
128'h000000000a3b29782578302c78257830, /* 2758 */
128'h782578302c302c7825287465736d656d, /* 2759 */
128'h464f5f4f4c43414d00000000000a3b29, /* 2760 */
128'h464f5f494843414d0000000054455346, /* 2761 */
128'h46464f5f524c50540000000054455346, /* 2762 */
128'h46464f5f534346540000000000544553, /* 2763 */
128'h4c5254434f49444d0000000000544553, /* 2764 */
128'h46464f5f534346520054455346464f5f, /* 2765 */
128'h5346464f5f5253520000000000544553, /* 2766 */
128'h46464f5f444142520000000000005445, /* 2767 */
128'h46464f5f524c50520000000000544553, /* 2768 */
128'h000000003f3f3f3f0000000000544553, /* 2769 */
128'h000064252b54455346464f5f524c5052, /* 2770 */
128'h6f746f72502050490000000000000047, /* 2771 */
128'h00000000000000000a50495049203d20, /* 2772 */
128'h6f746f72502050490000000000000054, /* 2773 */
128'h6f746f7250205049000a504745203d20, /* 2774 */
128'h6165682074736574000a505550203d20, /* 2775 */
128'h6e6f6320747365740000000a3a726564, /* 2776 */
128'h6f746f7250205049000a3a73746e6574, /* 2777 */
128'h6f746f7250205049000a504449203d20, /* 2778 */
128'h6f746f725020504900000a5054203d20, /* 2779 */
128'h00000000000000000a50434344203d20, /* 2780 */
128'h6f746f72502050490000000000000036, /* 2781 */
128'h00000000000000000a50565352203d20, /* 2782 */
128'h000a455247203d206f746f7250205049, /* 2783 */
128'h000a505345203d206f746f7250205049, /* 2784 */
128'h00000a4841203d206f746f7250205049, /* 2785 */
128'h000a50544d203d206f746f7250205049, /* 2786 */
128'h5054454542203d206f746f7250205049, /* 2787 */
128'h6f746f72502050490000000000000a48, /* 2788 */
128'h000000000000000a5041434e45203d20, /* 2789 */
128'h6f746f7250205049000000000000004d, /* 2790 */
128'h00000000000000000a504d4f43203d20, /* 2791 */
128'h0a50544353203d206f746f7250205049, /* 2792 */
128'h6f746f72502050490000000000000000, /* 2793 */
128'h00000000000a4554494c504455203d20, /* 2794 */
128'h0a534c504d203d206f746f7250205049, /* 2795 */
128'h6f746f72502050490000000000000000, /* 2796 */
128'h6f746f7270205049000a574152203d20, /* 2797 */
128'h2820646574726f707075736e75203d20, /* 2798 */
128'h79745f6f746f7270000000000a297825, /* 2799 */
128'h0000000000000a78257830203d206570, /* 2800 */
128'h727265746e692064656c646e61686e75, /* 2801 */
128'h414d2070757465530000000a21747075, /* 2802 */
128'h4d454f2049505351000a726464612043, /* 2803 */
128'h0000000000000a7825203d205d64255b, /* 2804 */
128'h00000a786c253a786c25203d2043414d, /* 2805 */
128'h3025203d20737365726464612043414d, /* 2806 */
128'h3230253a783230253a783230253a7832, /* 2807 */
128'h0000000a2e783230253a783230253a78, /* 2808 */
128'h00007f7c5d5b3f3e3d3c3b3a2c2b2a22, /* 2809 */
128'h007f7c5d5b3f3e3d3c3b3a2e2c2b2a22, /* 2810 */
128'h66656463626139383736353433323130, /* 2811 */
128'h72776f6c2f6372730000000000000000, /* 2812 */
128'h00000000000000632e636d6d5f637369, /* 2813 */
128'h61625f6473203d3d20657361625f6473, /* 2814 */
128'h5f63736972776f6c00726464615f6573, /* 2815 */
128'h000a74756f656d6974207325203a6473, /* 2816 */
128'h616d202c6465766f6d65722064726143, /* 2817 */
128'h6425206f74206465676e616863206b73, /* 2818 */
128'h736e692064726143000000000000000a, /* 2819 */
128'h6e616863206b73616d202c6465747265, /* 2820 */
128'h0000000000000a6425206f7420646567, /* 2821 */
128'h25207461206465746165726320636d6d, /* 2822 */
128'h0000000a7825203d2074736f68202c78, /* 2823 */
128'h0000000000006f4e0000000000736559, /* 2824 */
128'h002020203a434d4d0000000052444420, /* 2825 */
128'h00000000000a7325203a656369766544, /* 2826 */
128'h3a4449207265727574636166756e614d, /* 2827 */
128'h0a7825203a4d454f000000000a782520, /* 2828 */
128'h6325203a656d614e0000000000000000, /* 2829 */
128'h0000000000000a206325632563256325, /* 2830 */
128'h00000a6425203a646565705320737542, /* 2831 */
128'h25203a79746963617061432068676948, /* 2832 */
128'h79746963617061430000000000000a73, /* 2833 */
128'h7464695720737542000000000000203a, /* 2834 */
128'h000000000a73257469622d6425203a68, /* 2835 */
128'h0000007825782520000000203a78250a, /* 2836 */
128'h00000000000064735f63736972776f6c, /* 2837 */
128'h0000000065646f6d206e776f6e6b6e55, /* 2838 */
128'h7830203a726f72724520737574617453, /* 2839 */
128'h2074756f656d69540000000a58383025, /* 2840 */
128'h616572206472616320676e6974696177, /* 2841 */
128'h6c69616620636d6d00000000000a7964, /* 2842 */
128'h6d6320706f747320646e6573206f7420, /* 2843 */
128'h6f6c62203a434d4d0000000000000a64, /* 2844 */
128'h20786c257830207265626d756e206b63, /* 2845 */
128'h6c2578302878616d2073646565637865, /* 2846 */
128'h203d3e20434d4d6500000000000a2978, /* 2847 */
128'h726f6620646572697571657220342e34, /* 2848 */
128'h642072657375206465636e61686e6520, /* 2849 */
128'h000000000000000a6165726120617461, /* 2850 */
128'h757320746f6e2073656f642064726143, /* 2851 */
128'h696e6f697469747261702074726f7070, /* 2852 */
128'h656f64206472614300000000000a676e, /* 2853 */
128'h20434820656e6966656420746f6e2073, /* 2854 */
128'h00000a657a69732070756f7267205057, /* 2855 */
128'h636e61686e6520617461642072657355, /* 2856 */
128'h5720434820746f6e2061657261206465, /* 2857 */
128'h696c6120657a69732070756f72672050, /* 2858 */
128'h72617020692550470000000a64656e67, /* 2859 */
128'h505720434820746f6e206e6f69746974, /* 2860 */
128'h67696c6120657a69732070756f726720, /* 2861 */
128'h656f642064726143000000000a64656e, /* 2862 */
128'h6e652074726f7070757320746f6e2073, /* 2863 */
128'h657475626972747461206465636e6168, /* 2864 */
128'h6e65206c61746f54000000000000000a, /* 2865 */
128'h6563786520657a6973206465636e6168, /* 2866 */
128'h20752528206d756d6978616d20736465, /* 2867 */
128'h656f64206472614300000a297525203e, /* 2868 */
128'h6f682074726f7070757320746f6e2073, /* 2869 */
128'h61702064656c6c6f72746e6f63207473, /* 2870 */
128'h6572206574697277206e6f6974697472, /* 2871 */
128'h6e6974746573207974696c696261696c, /* 2872 */
128'h726c61206472614300000000000a7367, /* 2873 */
128'h64656e6f697469747261702079646165, /* 2874 */
128'h206f6e203a434d4d000000000000000a, /* 2875 */
128'h0000000a746e65736572702064726163, /* 2876 */
128'h73657220746f6e206469642064726143, /* 2877 */
128'h20656761746c6f76206f7420646e6f70, /* 2878 */
128'h00000000000000000a217463656c6573, /* 2879 */
128'h7463656c6573206f7420656c62616e75, /* 2880 */
128'h00000000000000000a65646f6d206120, /* 2881 */
128'h646e756f66206473635f747865206f4e, /* 2882 */
128'h78363025206e614d0000000000000a21, /* 2883 */
128'h000000783430257834302520726e5320, /* 2884 */
128'h00000000632563256325632563256325, /* 2885 */
128'h6167656c20434d4d00000064252e6425, /* 2886 */
128'h636167654c2044530000000000007963, /* 2887 */
128'h6867694820434d4d0000000000000079, /* 2888 */
128'h0000297a484d36322820646565705320, /* 2889 */
128'h35282064656570532068676948204453, /* 2890 */
128'h6867694820434d4d000000297a484d30, /* 2891 */
128'h0000297a484d32352820646565705320, /* 2892 */
128'h7a484d32352820323552444420434d4d, /* 2893 */
128'h31524453205348550000000000000029, /* 2894 */
128'h00000000000000297a484d3532282032, /* 2895 */
128'h7a484d30352820353252445320534855, /* 2896 */
128'h35524453205348550000000000000029, /* 2897 */
128'h000000000000297a484d303031282030, /* 2898 */
128'h7a484d30352820303552444420534855, /* 2899 */
128'h31524453205348550000000000000029, /* 2900 */
128'h0000000000297a484d38303228203430, /* 2901 */
128'h0000297a484d30303228203030325348, /* 2902 */
128'h6f6e2064252065636976654420434d4d, /* 2903 */
128'h00000000000000000a646e756f662074, /* 2904 */
128'h000000000000445300000000434d4d65, /* 2905 */
128'h000000297325282000006425203a7325, /* 2906 */
128'h6e656c20656c69460000000000636d6d, /* 2907 */
128'h000000000000000a6425203d20687467, /* 2908 */
128'h0a7325203d202964252c70252835646d, /* 2909 */
128'h666c652064616f6c0000000000000000, /* 2910 */
128'h000a79726f6d656d20524444206f7420, /* 2911 */
128'h2064656c696166206461657220666c65, /* 2912 */
128'h000000646c252065646f632068746977, /* 2913 */
128'h6f6f7420687461702074736575716552, /* 2914 */
128'h00000000000a646c25202e676e6f6c20, /* 2915 */
128'h732522203a717277000000000000002f, /* 2916 */
128'h0a64253d657a69736b636f6c62202c22, /* 2917 */
128'h20657669656365520000000000000000, /* 2918 */
128'h0000000000000a2e646e6520656c6966, /* 2919 */
128'h656c6c6163207172775f656c646e6168, /* 2920 */
128'h206c6167656c6c4900000000000a2e64, /* 2921 */
128'h0a2e6e6f6974617265706f2050544654, /* 2922 */
128'h75716572206e656c0000000000000000, /* 2923 */
128'h6175746361202c5825203d2064657269, /* 2924 */
128'h000000005c2d2f7c000a7825203d206c, /* 2925 */
128'h20646564616f6c2065687420746f6f42, /* 2926 */
128'h6572646461207461206d6172676f7270, /* 2927 */
128'h000000000000000a2e2e2e7025207373, /* 2928 */
128'h445320746e756f6d206f74206c696146, /* 2929 */
128'h000000000000000a2172657669726420, /* 2930 */
128'h6e69206e69622e746f6f622064616f4c, /* 2931 */
128'h0000000000000a79726f6d656d206f74, /* 2932 */
128'h00000000000000006e69622e746f6f62, /* 2933 */
128'h62206e65706f206f742064656c696146, /* 2934 */
128'h206f74206c6961660000000a21746f6f, /* 2935 */
128'h000000000021656c69662065736f6c63, /* 2936 */
128'h6420746e756f6d75206f74206c696166, /* 2937 */
128'h20746f6f622d750a00000000216b7369, /* 2938 */
128'h67617473207473726966206465736162, /* 2939 */
128'h00000a726564616f6c20746f6f622065, /* 2940 */
128'h696166207325206e6f69747265737361, /* 2941 */
128'h696c202c732520656c6966202c64656c, /* 2942 */
128'h206e6f6974636e7566202c642520656e, /* 2943 */
128'h3a4552554c49414600000000000a7325, /* 2944 */
128'h74612078257830203d21207825783020, /* 2945 */
128'h00000a2e782578302074657366666f20, /* 2946 */
128'h7025203d203270202c7025203d203170, /* 2947 */
128'h2020202020202020000000000000000a, /* 2948 */
128'h08080808080808080000000000202020, /* 2949 */
128'h20676e69747465730000000000080808, /* 2950 */
128'h20676e69747365740000000000007525, /* 2951 */
128'h3a4552554c4941460000000000007525, /* 2952 */
128'h64612064616220656c626973736f7020, /* 2953 */
128'h666f20746120656e696c207373657264, /* 2954 */
128'h00000000000a2e782578302074657366, /* 2955 */
128'h7478656e206f7420676e697070696b53, /* 2956 */
128'h000000000000000a2e2e2e7473657420, /* 2957 */
128'h20202020200808080808080808080808, /* 2958 */
128'h08080808080808080808202020202020, /* 2959 */
128'h00000000000820080000000000000008, /* 2960 */
128'h78302073692065676e61722074736574, /* 2961 */
128'h00000000000a70257830206f74207025, /* 2962 */
128'h000000000075252f00752520706f6f4c, /* 2963 */
128'h6441206b637574530000000000000a3a, /* 2964 */
128'h0000203a732520200000007373657264, /* 2965 */
128'h00000a2e656e6f4400000000000a6b6f, /* 2966 */
128'h4d415244206c6174656d20657261420a, /* 2967 */
128'h65747365746d656d00000a7473657420, /* 2968 */
128'h20302e332e34206e6f69737265762072, /* 2969 */
128'h000000000000000a297469622d642528, /* 2970 */
128'h30322029432820746867697279706f43, /* 2971 */
128'h2073656c7261684320323130322d3130, /* 2972 */
128'h000000000000000a2e6e6f62617a6143, /* 2973 */
128'h74207265646e75206465736e6563694c, /* 2974 */
128'h50206c6172656e654720554e47206568, /* 2975 */
128'h65762065736e6563694c2063696c6275, /* 2976 */
128'h0a2e29796c6e6f282032206e6f697372, /* 2977 */
128'h5f676e696b726f770000000000000000, /* 2978 */
128'h20646c25202c424b6425203d20746573, /* 2979 */
128'h6c25202c736e6f697463757274736e69, /* 2980 */
128'h203d20495043202c73656c6379632064, /* 2981 */
128'h00000000000000000a646c252e646c25, /* 2982 */
128'h46454443424139383736353433323130, /* 2983 */
128'h6f57206f6c6c65480000000000000000, /* 2984 */
128'h205d64255b70777300000a0d21646c72, /* 2985 */
128'h73206863746977530000000a5825203d, /* 2986 */
128'h000a58252c5825203d20676e69747465, /* 2987 */
128'h5825203d2064656573206d6f646e6152, /* 2988 */
128'h0a746f6f62204453000000000000000a, /* 2989 */
128'h6f6f6220495053510000000000000000, /* 2990 */
128'h736574204d4152440000000000000a74, /* 2991 */
128'h6f6f6220505446540000000000000a74, /* 2992 */
128'h65742065686361430000000000000a74, /* 2993 */
128'h00000a0d7061727400000000000a7473, /* 2994 */
128'h00000002464c457fcccccccccccccccd, /* 2995 */
128'h1032547698badcfeefcdab8967452301, /* 2996 */
128'h5851f42d4c957f2d1000000020000000, /* 2997 */
128'haaaaaaaaaaaaaaaa5555555555555555, /* 2998 */
128'h00000000000000000000000000000000, /* 2999 */
128'h00000000000000000000000000000000, /* 3000 */
128'h00000000000000000000000000000000, /* 3001 */
128'h00000000000000000000000000000000, /* 3002 */
128'h00000000000000000000000000000000, /* 3003 */
128'h00000000000000000000000000000000, /* 3004 */
128'h00000000000000000000000000000000, /* 3005 */
128'h00000000000000000000000000000000, /* 3006 */
128'h00000000000000000000000000000000, /* 3007 */
128'h00004b4d47545045000000030f060301, /* 3008 */
128'h000000004300000000000000004b4d47, /* 3009 */
128'h00000000ffffffff0000000000000000, /* 3010 */
128'h0000646d635f6473000000000c000000, /* 3011 */
128'h00000000ffffffff00006772615f6473, /* 3012 */
128'h000000002f7c5c2d0000000087feb3f8, /* 3013 */
128'h000000060000000087feb5b0cc33aa55, /* 3014 */
128'h87fe70980000000000000000ffffffff, /* 3015 */
128'h00000000000000000000000000000000, /* 3016 */
128'h00000000000000000000000000000000, /* 3017 */
128'h00000000000000000000000000000000, /* 3018 */
128'h00000000000000000000000000000000, /* 3019 */
128'h00000000000000000000000000000000, /* 3020 */
128'h00000000000000000000000000000000, /* 3021 */
128'h00000000000000000000000000000000, /* 3022 */
128'h00000000000000000000000000000000, /* 3023 */
128'h00000000000000000000000000000000, /* 3024 */
128'h00000000000000000000000000000000, /* 3025 */
128'h00000000000000000000000000000000, /* 3026 */
128'h00000000000000000000000000000000, /* 3027 */
128'h00000000000000000000000000000000, /* 3028 */
128'h00000000000000000000000000000000, /* 3029 */
128'h00000000000000000000000000000000, /* 3030 */
128'h00000000000000000000000000000000, /* 3031 */
128'h00000000000000000000000000000000, /* 3032 */
128'h00000000000000000000000000000000, /* 3033 */
128'h00000000000000000000000000000000, /* 3034 */
128'h00000000000000000000000000000000, /* 3035 */
128'h00000000000000000000000000000000, /* 3036 */
128'h00000000000000000000000000000000, /* 3037 */
128'h00000000000000000000000000000000, /* 3038 */
128'h00000000000000000000000000000000, /* 3039 */
128'h00000000000000000000000000000000, /* 3040 */
128'h00000000000000000000000000000000, /* 3041 */
128'h00000000000000000000000000000000, /* 3042 */
128'h00000000000000000000000000000000, /* 3043 */
128'h00000000000000000000000000000000, /* 3044 */
128'h00000000000000000000000000000000, /* 3045 */
128'h00000000000000000000000000000000, /* 3046 */
128'h00000000000000000000000000000000, /* 3047 */
128'h00000000000000000000000000000000, /* 3048 */
128'h00000000000000000000000000000000, /* 3049 */
128'h00000000000000000000000000000000, /* 3050 */
128'h00000000000000000000000000000000, /* 3051 */
128'h00000000000000000000000000000000, /* 3052 */
128'h00000000000000000000000000000000, /* 3053 */
128'h00000000000000000000000000000000, /* 3054 */
128'h00000000000000000000000000000000, /* 3055 */
128'h00000000000000000000000000000000, /* 3056 */
128'h00000000000000000000000000000000, /* 3057 */
128'h00000000000000000000000000000000, /* 3058 */
128'h00000000000000000000000000000000, /* 3059 */
128'h00000000000000000000000000000000, /* 3060 */
128'h00000000000000000000000000000000, /* 3061 */
128'h00000000000000000000000000000000, /* 3062 */
128'h00000000000000000000000000000000, /* 3063 */
128'h00000000000000000000000000000000, /* 3064 */
128'h00000000000000000000000000000000, /* 3065 */
128'h00000000000000000000000000000000, /* 3066 */
128'h00000000000000000000000000000000, /* 3067 */
128'h00000000000000000000000000000000, /* 3068 */
128'h00000000000000000000000000000000, /* 3069 */
128'h00000000000000000000000000000000, /* 3070 */
128'h00000000000000000000000000000000, /* 3071 */
128'h00000000000000000000000000000000, /* 3072 */
128'h00000000000000000000000000000000, /* 3073 */
128'h00000000000000000000000000000000, /* 3074 */
128'h00000000000000000000000000000000, /* 3075 */
128'h00000000000000000000000000000000, /* 3076 */
128'h00000000000000000000000000000000, /* 3077 */
128'h00000000000000000000000000000000, /* 3078 */
128'h00000000000000000000000000000000, /* 3079 */
128'h00000000000000000000000000000000, /* 3080 */
128'h00000000000000000000000000000000, /* 3081 */
128'h00000000000000000000000000000000, /* 3082 */
128'h00000000000000000000000000000000, /* 3083 */
128'h00000000000000000000000000000000, /* 3084 */
128'h00000000000000000000000000000000, /* 3085 */
128'h00000000000000000000000000000000, /* 3086 */
128'h00000000000000000000000000000000, /* 3087 */
128'h00000000000000000000000000000000, /* 3088 */
128'h00000000000000000000000000000000, /* 3089 */
128'h00000000000000000000000000000000, /* 3090 */
128'h00000000000000000000000000000000, /* 3091 */
128'h00000000000000000000000000000000, /* 3092 */
128'h00000000000000000000000000000000, /* 3093 */
128'h00000000000000000000000000000000, /* 3094 */
128'h00000000000000000000000000000000, /* 3095 */
128'h00000000000000000000000000000000, /* 3096 */
128'h00000000000000000000000000000000, /* 3097 */
128'h00000000000000000000000000000000, /* 3098 */
128'h00000000000000000000000000000000, /* 3099 */
128'h00000000000000000000000000000000, /* 3100 */
128'h00000000000000000000000000000000, /* 3101 */
128'h00000000000000000000000000000000, /* 3102 */
128'h00000000000000000000000000000000, /* 3103 */
128'h00000000000000000000000000000000, /* 3104 */
128'h00000000000000000000000000000000, /* 3105 */
128'h00000000000000000000000000000000, /* 3106 */
128'h00000000000000000000000000000000, /* 3107 */
128'h00000000000000000000000000000000, /* 3108 */
128'h00000000000000000000000000000000, /* 3109 */
128'h00000000000000000000000000000000, /* 3110 */
128'h00000000000000000000000000000000, /* 3111 */
128'h00000000000000000000000000000000, /* 3112 */
128'h00000000000000000000000000000000, /* 3113 */
128'h00000000000000000000000000000000, /* 3114 */
128'h00000000000000000000000000000000, /* 3115 */
128'h00000000000000000000000000000000, /* 3116 */
128'h00000000000000000000000000000000, /* 3117 */
128'h00000000000000000000000000000000, /* 3118 */
128'h00000000000000000000000000000000, /* 3119 */
128'h00000000000000000000000000000000, /* 3120 */
128'h00000000000000000000000000000000, /* 3121 */
128'h00000000000000000000000000000000, /* 3122 */
128'h00000000000000000000000000000000, /* 3123 */
128'h00000000000000000000000000000000, /* 3124 */
128'h00000000000000000000000000000000, /* 3125 */
128'h00000000000000000000000000000000, /* 3126 */
128'h00000000000000000000000000000000, /* 3127 */
128'h00000000000000000000000000000000, /* 3128 */
128'h00000000000000000000000000000000, /* 3129 */
128'h00000000000000000000000000000000, /* 3130 */
128'h00000000000000000000000000000000, /* 3131 */
128'h00000000000000000000000000000000, /* 3132 */
128'h00000000000000000000000000000000, /* 3133 */
128'h00000000000000000000000000000000, /* 3134 */
128'h00000000000000000000000000000000, /* 3135 */
128'h00000000000000000000000000000000, /* 3136 */
128'h00000000000000000000000000000000, /* 3137 */
128'h00000000000000000000000000000000, /* 3138 */
128'h00000000000000000000000000000000, /* 3139 */
128'h00000000000000000000000000000000, /* 3140 */
128'h00000000000000000000000000000000, /* 3141 */
128'h00000000000000000000000000000000, /* 3142 */
128'h00000000000000000000000000000000, /* 3143 */
128'h00000000000000000000000000000000, /* 3144 */
128'h00000000000000000000000000000000, /* 3145 */
128'h00000000000000000000000000000000, /* 3146 */
128'h00000000000000000000000000000000, /* 3147 */
128'h00000000000000000000000000000000, /* 3148 */
128'h00000000000000000000000000000000, /* 3149 */
128'h00000000000000000000000000000000, /* 3150 */
128'h00000000000000000000000000000000, /* 3151 */
128'h00000000000000000000000000000000, /* 3152 */
128'h00000000000000000000000000000000, /* 3153 */
128'h00000000000000000000000000000000, /* 3154 */
128'h00000000000000000000000000000000, /* 3155 */
128'h00000000000000000000000000000000, /* 3156 */
128'h00000000000000000000000000000000, /* 3157 */
128'h00000000000000000000000000000000, /* 3158 */
128'h00000000000000000000000000000000, /* 3159 */
128'h00000000000000000000000000000000, /* 3160 */
128'h00000000000000000000000000000000, /* 3161 */
128'h00000000000000000000000000000000, /* 3162 */
128'h00000000000000000000000000000000, /* 3163 */
128'h00000000000000000000000000000000, /* 3164 */
128'h00000000000000000000000000000000, /* 3165 */
128'h00000000000000000000000000000000, /* 3166 */
128'h00000000000000000000000000000000, /* 3167 */
128'h00000000000000000000000000000000, /* 3168 */
128'h00000000000000000000000000000000, /* 3169 */
128'h00000000000000000000000000000000, /* 3170 */
128'h00000000000000000000000000000000, /* 3171 */
128'h00000000000000000000000000000000, /* 3172 */
128'h00000000000000000000000000000000, /* 3173 */
128'h00000000000000000000000000000000, /* 3174 */
128'h00000000000000000000000000000000, /* 3175 */
128'h00000000000000000000000000000000, /* 3176 */
128'h00000000000000000000000000000000, /* 3177 */
128'h00000000000000000000000000000000, /* 3178 */
128'h00000000000000000000000000000000, /* 3179 */
128'h00000000000000000000000000000000, /* 3180 */
128'h00000000000000000000000000000000, /* 3181 */
128'h00000000000000000000000000000000, /* 3182 */
128'h00000000000000000000000000000000, /* 3183 */
128'h00000000000000000000000000000000, /* 3184 */
128'h00000000000000000000000000000000, /* 3185 */
128'h00000000000000000000000000000000, /* 3186 */
128'h00000000000000000000000000000000, /* 3187 */
128'h00000000000000000000000000000000, /* 3188 */
128'h00000000000000000000000000000000, /* 3189 */
128'h00000000000000000000000000000000, /* 3190 */
128'h00000000000000000000000000000000, /* 3191 */
128'h00000000000000000000000000000000, /* 3192 */
128'h00000000000000000000000000000000, /* 3193 */
128'h00000000000000000000000000000000, /* 3194 */
128'h00000000000000000000000000000000, /* 3195 */
128'h00000000000000000000000000000000, /* 3196 */
128'h00000000000000000000000000000000, /* 3197 */
128'h00000000000000000000000000000000, /* 3198 */
128'h00000000000000000000000000000000, /* 3199 */
128'h00000000000000000000000000000000, /* 3200 */
128'h00000000000000000000000000000000, /* 3201 */
128'h00000000000000000000000000000000, /* 3202 */
128'h00000000000000000000000000000000, /* 3203 */
128'h00000000000000000000000000000000, /* 3204 */
128'h00000000000000000000000000000000, /* 3205 */
128'h00000000000000000000000000000000, /* 3206 */
128'h00000000000000000000000000000000, /* 3207 */
128'h00000000000000000000000000000000, /* 3208 */
128'h00000000000000000000000000000000, /* 3209 */
128'h00000000000000000000000000000000, /* 3210 */
128'h00000000000000000000000000000000, /* 3211 */
128'h00000000000000000000000000000000, /* 3212 */
128'h00000000000000000000000000000000, /* 3213 */
128'h00000000000000000000000000000000, /* 3214 */
128'h00000000000000000000000000000000, /* 3215 */
128'h00000000000000000000000000000000, /* 3216 */
128'h00000000000000000000000000000000, /* 3217 */
128'h00000000000000000000000000000000, /* 3218 */
128'h00000000000000000000000000000000, /* 3219 */
128'h00000000000000000000000000000000, /* 3220 */
128'h00000000000000000000000000000000, /* 3221 */
128'h00000000000000000000000000000000, /* 3222 */
128'h00000000000000000000000000000000, /* 3223 */
128'h00000000000000000000000000000000, /* 3224 */
128'h00000000000000000000000000000000, /* 3225 */
128'h00000000000000000000000000000000, /* 3226 */
128'h00000000000000000000000000000000, /* 3227 */
128'h00000000000000000000000000000000, /* 3228 */
128'h00000000000000000000000000000000, /* 3229 */
128'h00000000000000000000000000000000, /* 3230 */
128'h00000000000000000000000000000000, /* 3231 */
128'h00000000000000000000000000000000, /* 3232 */
128'h00000000000000000000000000000000, /* 3233 */
128'h00000000000000000000000000000000, /* 3234 */
128'h00000000000000000000000000000000, /* 3235 */
128'h00000000000000000000000000000000, /* 3236 */
128'h00000000000000000000000000000000, /* 3237 */
128'h00000000000000000000000000000000, /* 3238 */
128'h00000000000000000000000000000000, /* 3239 */
128'h00000000000000000000000000000000, /* 3240 */
128'h00000000000000000000000000000000, /* 3241 */
128'h00000000000000000000000000000000, /* 3242 */
128'h00000000000000000000000000000000, /* 3243 */
128'h00000000000000000000000000000000, /* 3244 */
128'h00000000000000000000000000000000, /* 3245 */
128'h00000000000000000000000000000000, /* 3246 */
128'h00000000000000000000000000000000, /* 3247 */
128'h00000000000000000000000000000000, /* 3248 */
128'h00000000000000000000000000000000, /* 3249 */
128'h00000000000000000000000000000000, /* 3250 */
128'h00000000000000000000000000000000, /* 3251 */
128'h00000000000000000000000000000000, /* 3252 */
128'h00000000000000000000000000000000, /* 3253 */
128'h00000000000000000000000000000000, /* 3254 */
128'h00000000000000000000000000000000, /* 3255 */
128'h00000000000000000000000000000000, /* 3256 */
128'h00000000000000000000000000000000, /* 3257 */
128'h00000000000000000000000000000000, /* 3258 */
128'h00000000000000000000000000000000, /* 3259 */
128'h00000000000000000000000000000000, /* 3260 */
128'h00000000000000000000000000000000, /* 3261 */
128'h00000000000000000000000000000000, /* 3262 */
128'h00000000000000000000000000000000, /* 3263 */
128'h00000000000000000000000000000000, /* 3264 */
128'h00000000000000000000000000000000, /* 3265 */
128'h00000000000000000000000000000000, /* 3266 */
128'h00000000000000000000000000000000, /* 3267 */
128'h00000000000000000000000000000000, /* 3268 */
128'h00000000000000000000000000000000, /* 3269 */
128'h00000000000000000000000000000000, /* 3270 */
128'h00000000000000000000000000000000, /* 3271 */
128'h00000000000000000000000000000000, /* 3272 */
128'h00000000000000000000000000000000, /* 3273 */
128'h00000000000000000000000000000000, /* 3274 */
128'h00000000000000000000000000000000, /* 3275 */
128'h00000000000000000000000000000000, /* 3276 */
128'h00000000000000000000000000000000, /* 3277 */
128'h00000000000000000000000000000000, /* 3278 */
128'h00000000000000000000000000000000, /* 3279 */
128'h00000000000000000000000000000000, /* 3280 */
128'h00000000000000000000000000000000, /* 3281 */
128'h00000000000000000000000000000000, /* 3282 */
128'h00000000000000000000000000000000, /* 3283 */
128'h00000000000000000000000000000000, /* 3284 */
128'h00000000000000000000000000000000, /* 3285 */
128'h00000000000000000000000000000000, /* 3286 */
128'h00000000000000000000000000000000, /* 3287 */
128'h00000000000000000000000000000000, /* 3288 */
128'h00000000000000000000000000000000, /* 3289 */
128'h00000000000000000000000000000000, /* 3290 */
128'h00000000000000000000000000000000, /* 3291 */
128'h00000000000000000000000000000000, /* 3292 */
128'h00000000000000000000000000000000, /* 3293 */
128'h00000000000000000000000000000000, /* 3294 */
128'h00000000000000000000000000000000, /* 3295 */
128'h00000000000000000000000000000000, /* 3296 */
128'h00000000000000000000000000000000, /* 3297 */
128'h00000000000000000000000000000000, /* 3298 */
128'h00000000000000000000000000000000, /* 3299 */
128'h00000000000000000000000000000000, /* 3300 */
128'h00000000000000000000000000000000, /* 3301 */
128'h00000000000000000000000000000000, /* 3302 */
128'h00000000000000000000000000000000, /* 3303 */
128'h00000000000000000000000000000000, /* 3304 */
128'h00000000000000000000000000000000, /* 3305 */
128'h00000000000000000000000000000000, /* 3306 */
128'h00000000000000000000000000000000, /* 3307 */
128'h00000000000000000000000000000000, /* 3308 */
128'h00000000000000000000000000000000, /* 3309 */
128'h00000000000000000000000000000000, /* 3310 */
128'h00000000000000000000000000000000, /* 3311 */
128'h00000000000000000000000000000000, /* 3312 */
128'h00000000000000000000000000000000, /* 3313 */
128'h00000000000000000000000000000000, /* 3314 */
128'h00000000000000000000000000000000, /* 3315 */
128'h00000000000000000000000000000000, /* 3316 */
128'h00000000000000000000000000000000, /* 3317 */
128'h00000000000000000000000000000000, /* 3318 */
128'h00000000000000000000000000000000, /* 3319 */
128'h00000000000000000000000000000000, /* 3320 */
128'h00000000000000000000000000000000, /* 3321 */
128'h00000000000000000000000000000000, /* 3322 */
128'h00000000000000000000000000000000, /* 3323 */
128'h00000000000000000000000000000000, /* 3324 */
128'h00000000000000000000000000000000, /* 3325 */
128'h00000000000000000000000000000000, /* 3326 */
128'h00000000000000000000000000000000, /* 3327 */
128'h00000000000000000000000000000000, /* 3328 */
128'h00000000000000000000000000000000, /* 3329 */
128'h00000000000000000000000000000000, /* 3330 */
128'h00000000000000000000000000000000, /* 3331 */
128'h00000000000000000000000000000000, /* 3332 */
128'h00000000000000000000000000000000, /* 3333 */
128'h00000000000000000000000000000000, /* 3334 */
128'h00000000000000000000000000000000, /* 3335 */
128'h00000000000000000000000000000000, /* 3336 */
128'h00000000000000000000000000000000, /* 3337 */
128'h00000000000000000000000000000000, /* 3338 */
128'h00000000000000000000000000000000, /* 3339 */
128'h00000000000000000000000000000000, /* 3340 */
128'h00000000000000000000000000000000, /* 3341 */
128'h00000000000000000000000000000000, /* 3342 */
128'h00000000000000000000000000000000, /* 3343 */
128'h00000000000000000000000000000000, /* 3344 */
128'h00000000000000000000000000000000, /* 3345 */
128'h00000000000000000000000000000000, /* 3346 */
128'h00000000000000000000000000000000, /* 3347 */
128'h00000000000000000000000000000000, /* 3348 */
128'h00000000000000000000000000000000, /* 3349 */
128'h00000000000000000000000000000000, /* 3350 */
128'h00000000000000000000000000000000, /* 3351 */
128'h00000000000000000000000000000000, /* 3352 */
128'h00000000000000000000000000000000, /* 3353 */
128'h00000000000000000000000000000000, /* 3354 */
128'h00000000000000000000000000000000, /* 3355 */
128'h00000000000000000000000000000000, /* 3356 */
128'h00000000000000000000000000000000, /* 3357 */
128'h00000000000000000000000000000000, /* 3358 */
128'h00000000000000000000000000000000, /* 3359 */
128'h00000000000000000000000000000000, /* 3360 */
128'h00000000000000000000000000000000, /* 3361 */
128'h00000000000000000000000000000000, /* 3362 */
128'h00000000000000000000000000000000, /* 3363 */
128'h00000000000000000000000000000000, /* 3364 */
128'h00000000000000000000000000000000, /* 3365 */
128'h00000000000000000000000000000000, /* 3366 */
128'h00000000000000000000000000000000, /* 3367 */
128'h00000000000000000000000000000000, /* 3368 */
128'h00000000000000000000000000000000, /* 3369 */
128'h00000000000000000000000000000000, /* 3370 */
128'h00000000000000000000000000000000, /* 3371 */
128'h00000000000000000000000000000000, /* 3372 */
128'h00000000000000000000000000000000, /* 3373 */
128'h00000000000000000000000000000000, /* 3374 */
128'h00000000000000000000000000000000, /* 3375 */
128'h00000000000000000000000000000000, /* 3376 */
128'h00000000000000000000000000000000, /* 3377 */
128'h00000000000000000000000000000000, /* 3378 */
128'h00000000000000000000000000000000, /* 3379 */
128'h00000000000000000000000000000000, /* 3380 */
128'h00000000000000000000000000000000, /* 3381 */
128'h00000000000000000000000000000000, /* 3382 */
128'h00000000000000000000000000000000, /* 3383 */
128'h00000000000000000000000000000000, /* 3384 */
128'h00000000000000000000000000000000, /* 3385 */
128'h00000000000000000000000000000000, /* 3386 */
128'h00000000000000000000000000000000, /* 3387 */
128'h00000000000000000000000000000000, /* 3388 */
128'h00000000000000000000000000000000, /* 3389 */
128'h00000000000000000000000000000000, /* 3390 */
128'h00000000000000000000000000000000, /* 3391 */
128'h00000000000000000000000000000000, /* 3392 */
128'h00000000000000000000000000000000, /* 3393 */
128'h00000000000000000000000000000000, /* 3394 */
128'h00000000000000000000000000000000, /* 3395 */
128'h00000000000000000000000000000000, /* 3396 */
128'h00000000000000000000000000000000, /* 3397 */
128'h00000000000000000000000000000000, /* 3398 */
128'h00000000000000000000000000000000, /* 3399 */
128'h00000000000000000000000000000000, /* 3400 */
128'h00000000000000000000000000000000, /* 3401 */
128'h00000000000000000000000000000000, /* 3402 */
128'h00000000000000000000000000000000, /* 3403 */
128'h00000000000000000000000000000000, /* 3404 */
128'h00000000000000000000000000000000, /* 3405 */
128'h00000000000000000000000000000000, /* 3406 */
128'h00000000000000000000000000000000, /* 3407 */
128'h00000000000000000000000000000000, /* 3408 */
128'h00000000000000000000000000000000, /* 3409 */
128'h00000000000000000000000000000000, /* 3410 */
128'h00000000000000000000000000000000, /* 3411 */
128'h00000000000000000000000000000000, /* 3412 */
128'h00000000000000000000000000000000, /* 3413 */
128'h00000000000000000000000000000000, /* 3414 */
128'h00000000000000000000000000000000, /* 3415 */
128'h00000000000000000000000000000000, /* 3416 */
128'h00000000000000000000000000000000, /* 3417 */
128'h00000000000000000000000000000000, /* 3418 */
128'h00000000000000000000000000000000, /* 3419 */
128'h00000000000000000000000000000000, /* 3420 */
128'h00000000000000000000000000000000, /* 3421 */
128'h00000000000000000000000000000000, /* 3422 */
128'h00000000000000000000000000000000, /* 3423 */
128'h00000000000000000000000000000000, /* 3424 */
128'h00000000000000000000000000000000, /* 3425 */
128'h00000000000000000000000000000000, /* 3426 */
128'h00000000000000000000000000000000, /* 3427 */
128'h00000000000000000000000000000000, /* 3428 */
128'h00000000000000000000000000000000, /* 3429 */
128'h00000000000000000000000000000000, /* 3430 */
128'h00000000000000000000000000000000, /* 3431 */
128'h00000000000000000000000000000000, /* 3432 */
128'h00000000000000000000000000000000, /* 3433 */
128'h00000000000000000000000000000000, /* 3434 */
128'h00000000000000000000000000000000, /* 3435 */
128'h00000000000000000000000000000000, /* 3436 */
128'h00000000000000000000000000000000, /* 3437 */
128'h00000000000000000000000000000000, /* 3438 */
128'h00000000000000000000000000000000, /* 3439 */
128'h00000000000000000000000000000000, /* 3440 */
128'h00000000000000000000000000000000, /* 3441 */
128'h00000000000000000000000000000000, /* 3442 */
128'h00000000000000000000000000000000, /* 3443 */
128'h00000000000000000000000000000000, /* 3444 */
128'h00000000000000000000000000000000, /* 3445 */
128'h00000000000000000000000000000000, /* 3446 */
128'h00000000000000000000000000000000, /* 3447 */
128'h00000000000000000000000000000000, /* 3448 */
128'h00000000000000000000000000000000, /* 3449 */
128'h00000000000000000000000000000000, /* 3450 */
128'h00000000000000000000000000000000, /* 3451 */
128'h00000000000000000000000000000000, /* 3452 */
128'h00000000000000000000000000000000, /* 3453 */
128'h00000000000000000000000000000000, /* 3454 */
128'h00000000000000000000000000000000, /* 3455 */
128'h00000000000000000000000000000000, /* 3456 */
128'h00000000000000000000000000000000, /* 3457 */
128'h00000000000000000000000000000000, /* 3458 */
128'h00000000000000000000000000000000, /* 3459 */
128'h00000000000000000000000000000000, /* 3460 */
128'h00000000000000000000000000000000, /* 3461 */
128'h00000000000000000000000000000000, /* 3462 */
128'h00000000000000000000000000000000, /* 3463 */
128'h00000000000000000000000000000000, /* 3464 */
128'h00000000000000000000000000000000, /* 3465 */
128'h00000000000000000000000000000000, /* 3466 */
128'h00000000000000000000000000000000, /* 3467 */
128'h00000000000000000000000000000000, /* 3468 */
128'h00000000000000000000000000000000, /* 3469 */
128'h00000000000000000000000000000000, /* 3470 */
128'h00000000000000000000000000000000, /* 3471 */
128'h00000000000000000000000000000000, /* 3472 */
128'h00000000000000000000000000000000, /* 3473 */
128'h00000000000000000000000000000000, /* 3474 */
128'h00000000000000000000000000000000, /* 3475 */
128'h00000000000000000000000000000000, /* 3476 */
128'h00000000000000000000000000000000, /* 3477 */
128'h00000000000000000000000000000000, /* 3478 */
128'h00000000000000000000000000000000, /* 3479 */
128'h00000000000000000000000000000000, /* 3480 */
128'h00000000000000000000000000000000, /* 3481 */
128'h00000000000000000000000000000000, /* 3482 */
128'h00000000000000000000000000000000, /* 3483 */
128'h00000000000000000000000000000000, /* 3484 */
128'h00000000000000000000000000000000, /* 3485 */
128'h00000000000000000000000000000000, /* 3486 */
128'h00000000000000000000000000000000, /* 3487 */
128'h00000000000000000000000000000000, /* 3488 */
128'h00000000000000000000000000000000, /* 3489 */
128'h00000000000000000000000000000000, /* 3490 */
128'h00000000000000000000000000000000, /* 3491 */
128'h00000000000000000000000000000000, /* 3492 */
128'h00000000000000000000000000000000, /* 3493 */
128'h00000000000000000000000000000000, /* 3494 */
128'h00000000000000000000000000000000, /* 3495 */
128'h00000000000000000000000000000000, /* 3496 */
128'h00000000000000000000000000000000, /* 3497 */
128'h00000000000000000000000000000000, /* 3498 */
128'h00000000000000000000000000000000, /* 3499 */
128'h00000000000000000000000000000000, /* 3500 */
128'h00000000000000000000000000000000, /* 3501 */
128'h00000000000000000000000000000000, /* 3502 */
128'h00000000000000000000000000000000, /* 3503 */
128'h00000000000000000000000000000000, /* 3504 */
128'h00000000000000000000000000000000, /* 3505 */
128'h00000000000000000000000000000000, /* 3506 */
128'h00000000000000000000000000000000, /* 3507 */
128'h00000000000000000000000000000000, /* 3508 */
128'h00000000000000000000000000000000, /* 3509 */
128'h00000000000000000000000000000000, /* 3510 */
128'h00000000000000000000000000000000, /* 3511 */
128'h00000000000000000000000000000000, /* 3512 */
128'h00000000000000000000000000000000, /* 3513 */
128'h00000000000000000000000000000000, /* 3514 */
128'h00000000000000000000000000000000, /* 3515 */
128'h00000000000000000000000000000000, /* 3516 */
128'h00000000000000000000000000000000, /* 3517 */
128'h00000000000000000000000000000000, /* 3518 */
128'h00000000000000000000000000000000, /* 3519 */
128'h00000000000000000000000000000000, /* 3520 */
128'h00000000000000000000000000000000, /* 3521 */
128'h00000000000000000000000000000000, /* 3522 */
128'h00000000000000000000000000000000, /* 3523 */
128'h00000000000000000000000000000000, /* 3524 */
128'h00000000000000000000000000000000, /* 3525 */
128'h00000000000000000000000000000000, /* 3526 */
128'h00000000000000000000000000000000, /* 3527 */
128'h00000000000000000000000000000000, /* 3528 */
128'h00000000000000000000000000000000, /* 3529 */
128'h00000000000000000000000000000000, /* 3530 */
128'h00000000000000000000000000000000, /* 3531 */
128'h00000000000000000000000000000000, /* 3532 */
128'h00000000000000000000000000000000, /* 3533 */
128'h00000000000000000000000000000000, /* 3534 */
128'h00000000000000000000000000000000, /* 3535 */
128'h00000000000000000000000000000000, /* 3536 */
128'h00000000000000000000000000000000, /* 3537 */
128'h00000000000000000000000000000000, /* 3538 */
128'h00000000000000000000000000000000, /* 3539 */
128'h00000000000000000000000000000000, /* 3540 */
128'h00000000000000000000000000000000, /* 3541 */
128'h00000000000000000000000000000000, /* 3542 */
128'h00000000000000000000000000000000, /* 3543 */
128'h00000000000000000000000000000000, /* 3544 */
128'h00000000000000000000000000000000, /* 3545 */
128'h00000000000000000000000000000000, /* 3546 */
128'h00000000000000000000000000000000, /* 3547 */
128'h00000000000000000000000000000000, /* 3548 */
128'h00000000000000000000000000000000, /* 3549 */
128'h00000000000000000000000000000000, /* 3550 */
128'h00000000000000000000000000000000, /* 3551 */
128'h00000000000000000000000000000000, /* 3552 */
128'h00000000000000000000000000000000, /* 3553 */
128'h00000000000000000000000000000000, /* 3554 */
128'h00000000000000000000000000000000, /* 3555 */
128'h00000000000000000000000000000000, /* 3556 */
128'h00000000000000000000000000000000, /* 3557 */
128'h00000000000000000000000000000000, /* 3558 */
128'h00000000000000000000000000000000, /* 3559 */
128'h00000000000000000000000000000000, /* 3560 */
128'h00000000000000000000000000000000, /* 3561 */
128'h00000000000000000000000000000000, /* 3562 */
128'h00000000000000000000000000000000, /* 3563 */
128'h00000000000000000000000000000000, /* 3564 */
128'h00000000000000000000000000000000, /* 3565 */
128'h00000000000000000000000000000000, /* 3566 */
128'h00000000000000000000000000000000, /* 3567 */
128'h00000000000000000000000000000000, /* 3568 */
128'h00000000000000000000000000000000, /* 3569 */
128'h00000000000000000000000000000000, /* 3570 */
128'h00000000000000000000000000000000, /* 3571 */
128'h00000000000000000000000000000000, /* 3572 */
128'h00000000000000000000000000000000, /* 3573 */
128'h00000000000000000000000000000000, /* 3574 */
128'h00000000000000000000000000000000, /* 3575 */
128'h00000000000000000000000000000000, /* 3576 */
128'h00000000000000000000000000000000, /* 3577 */
128'h00000000000000000000000000000000, /* 3578 */
128'h00000000000000000000000000000000, /* 3579 */
128'h00000000000000000000000000000000, /* 3580 */
128'h00000000000000000000000000000000, /* 3581 */
128'h00000000000000000000000000000000, /* 3582 */
128'h00000000000000000000000000000000, /* 3583 */
128'h00000000000000000000000000000000, /* 3584 */
128'h00000000000000000000000000000000, /* 3585 */
128'h00000000000000000000000000000000, /* 3586 */
128'h00000000000000000000000000000000, /* 3587 */
128'h00000000000000000000000000000000, /* 3588 */
128'h00000000000000000000000000000000, /* 3589 */
128'h00000000000000000000000000000000, /* 3590 */
128'h00000000000000000000000000000000, /* 3591 */
128'h00000000000000000000000000000000, /* 3592 */
128'h00000000000000000000000000000000, /* 3593 */
128'h00000000000000000000000000000000, /* 3594 */
128'h00000000000000000000000000000000, /* 3595 */
128'h00000000000000000000000000000000, /* 3596 */
128'h00000000000000000000000000000000, /* 3597 */
128'h00000000000000000000000000000000, /* 3598 */
128'h00000000000000000000000000000000, /* 3599 */
128'h00000000000000000000000000000000, /* 3600 */
128'h00000000000000000000000000000000, /* 3601 */
128'h00000000000000000000000000000000, /* 3602 */
128'h00000000000000000000000000000000, /* 3603 */
128'h00000000000000000000000000000000, /* 3604 */
128'h00000000000000000000000000000000, /* 3605 */
128'h00000000000000000000000000000000, /* 3606 */
128'h00000000000000000000000000000000, /* 3607 */
128'h00000000000000000000000000000000, /* 3608 */
128'h00000000000000000000000000000000, /* 3609 */
128'h00000000000000000000000000000000, /* 3610 */
128'h00000000000000000000000000000000, /* 3611 */
128'h00000000000000000000000000000000, /* 3612 */
128'h00000000000000000000000000000000, /* 3613 */
128'h00000000000000000000000000000000, /* 3614 */
128'h00000000000000000000000000000000, /* 3615 */
128'h00000000000000000000000000000000, /* 3616 */
128'h00000000000000000000000000000000, /* 3617 */
128'h00000000000000000000000000000000, /* 3618 */
128'h00000000000000000000000000000000, /* 3619 */
128'h00000000000000000000000000000000, /* 3620 */
128'h00000000000000000000000000000000, /* 3621 */
128'h00000000000000000000000000000000, /* 3622 */
128'h00000000000000000000000000000000, /* 3623 */
128'h00000000000000000000000000000000, /* 3624 */
128'h00000000000000000000000000000000, /* 3625 */
128'h00000000000000000000000000000000, /* 3626 */
128'h00000000000000000000000000000000, /* 3627 */
128'h00000000000000000000000000000000, /* 3628 */
128'h00000000000000000000000000000000, /* 3629 */
128'h00000000000000000000000000000000, /* 3630 */
128'h00000000000000000000000000000000, /* 3631 */
128'h00000000000000000000000000000000, /* 3632 */
128'h00000000000000000000000000000000, /* 3633 */
128'h00000000000000000000000000000000, /* 3634 */
128'h00000000000000000000000000000000, /* 3635 */
128'h00000000000000000000000000000000, /* 3636 */
128'h00000000000000000000000000000000, /* 3637 */
128'h00000000000000000000000000000000, /* 3638 */
128'h00000000000000000000000000000000, /* 3639 */
128'h00000000000000000000000000000000, /* 3640 */
128'h00000000000000000000000000000000, /* 3641 */
128'h00000000000000000000000000000000, /* 3642 */
128'h00000000000000000000000000000000, /* 3643 */
128'h00000000000000000000000000000000, /* 3644 */
128'h00000000000000000000000000000000, /* 3645 */
128'h00000000000000000000000000000000, /* 3646 */
128'h00000000000000000000000000000000, /* 3647 */
128'h00000000000000000000000000000000, /* 3648 */
128'h00000000000000000000000000000000, /* 3649 */
128'h00000000000000000000000000000000, /* 3650 */
128'h00000000000000000000000000000000, /* 3651 */
128'h00000000000000000000000000000000, /* 3652 */
128'h00000000000000000000000000000000, /* 3653 */
128'h00000000000000000000000000000000, /* 3654 */
128'h00000000000000000000000000000000, /* 3655 */
128'h00000000000000000000000000000000, /* 3656 */
128'h00000000000000000000000000000000, /* 3657 */
128'h00000000000000000000000000000000, /* 3658 */
128'h00000000000000000000000000000000, /* 3659 */
128'h00000000000000000000000000000000, /* 3660 */
128'h00000000000000000000000000000000, /* 3661 */
128'h00000000000000000000000000000000, /* 3662 */
128'h00000000000000000000000000000000, /* 3663 */
128'h00000000000000000000000000000000, /* 3664 */
128'h00000000000000000000000000000000, /* 3665 */
128'h00000000000000000000000000000000, /* 3666 */
128'h00000000000000000000000000000000, /* 3667 */
128'h00000000000000000000000000000000, /* 3668 */
128'h00000000000000000000000000000000, /* 3669 */
128'h00000000000000000000000000000000, /* 3670 */
128'h00000000000000000000000000000000, /* 3671 */
128'h00000000000000000000000000000000, /* 3672 */
128'h00000000000000000000000000000000, /* 3673 */
128'h00000000000000000000000000000000, /* 3674 */
128'h00000000000000000000000000000000, /* 3675 */
128'h00000000000000000000000000000000, /* 3676 */
128'h00000000000000000000000000000000, /* 3677 */
128'h00000000000000000000000000000000, /* 3678 */
128'h00000000000000000000000000000000, /* 3679 */
128'h00000000000000000000000000000000, /* 3680 */
128'h00000000000000000000000000000000, /* 3681 */
128'h00000000000000000000000000000000, /* 3682 */
128'h00000000000000000000000000000000, /* 3683 */
128'h00000000000000000000000000000000, /* 3684 */
128'h00000000000000000000000000000000, /* 3685 */
128'h00000000000000000000000000000000, /* 3686 */
128'h00000000000000000000000000000000, /* 3687 */
128'h00000000000000000000000000000000, /* 3688 */
128'h00000000000000000000000000000000, /* 3689 */
128'h00000000000000000000000000000000, /* 3690 */
128'h00000000000000000000000000000000, /* 3691 */
128'h00000000000000000000000000000000, /* 3692 */
128'h00000000000000000000000000000000, /* 3693 */
128'h00000000000000000000000000000000, /* 3694 */
128'h00000000000000000000000000000000, /* 3695 */
128'h00000000000000000000000000000000, /* 3696 */
128'h00000000000000000000000000000000, /* 3697 */
128'h00000000000000000000000000000000, /* 3698 */
128'h00000000000000000000000000000000, /* 3699 */
128'h00000000000000000000000000000000, /* 3700 */
128'h00000000000000000000000000000000, /* 3701 */
128'h00000000000000000000000000000000, /* 3702 */
128'h00000000000000000000000000000000, /* 3703 */
128'h00000000000000000000000000000000, /* 3704 */
128'h00000000000000000000000000000000, /* 3705 */
128'h00000000000000000000000000000000, /* 3706 */
128'h00000000000000000000000000000000, /* 3707 */
128'h00000000000000000000000000000000, /* 3708 */
128'h00000000000000000000000000000000, /* 3709 */
128'h00000000000000000000000000000000, /* 3710 */
128'h00000000000000000000000000000000, /* 3711 */
128'h00000000000000000000000000000000, /* 3712 */
128'h00000000000000000000000000000000, /* 3713 */
128'h00000000000000000000000000000000, /* 3714 */
128'h00000000000000000000000000000000, /* 3715 */
128'h00000000000000000000000000000000, /* 3716 */
128'h00000000000000000000000000000000, /* 3717 */
128'h00000000000000000000000000000000, /* 3718 */
128'h00000000000000000000000000000000, /* 3719 */
128'h00000000000000000000000000000000, /* 3720 */
128'h00000000000000000000000000000000, /* 3721 */
128'h00000000000000000000000000000000, /* 3722 */
128'h00000000000000000000000000000000, /* 3723 */
128'h00000000000000000000000000000000, /* 3724 */
128'h00000000000000000000000000000000, /* 3725 */
128'h00000000000000000000000000000000, /* 3726 */
128'h00000000000000000000000000000000, /* 3727 */
128'h00000000000000000000000000000000, /* 3728 */
128'h00000000000000000000000000000000, /* 3729 */
128'h00000000000000000000000000000000, /* 3730 */
128'h00000000000000000000000000000000, /* 3731 */
128'h00000000000000000000000000000000, /* 3732 */
128'h00000000000000000000000000000000, /* 3733 */
128'h00000000000000000000000000000000, /* 3734 */
128'h00000000000000000000000000000000, /* 3735 */
128'h00000000000000000000000000000000, /* 3736 */
128'h00000000000000000000000000000000, /* 3737 */
128'h00000000000000000000000000000000, /* 3738 */
128'h00000000000000000000000000000000, /* 3739 */
128'h00000000000000000000000000000000, /* 3740 */
128'h00000000000000000000000000000000, /* 3741 */
128'h00000000000000000000000000000000, /* 3742 */
128'h00000000000000000000000000000000, /* 3743 */
128'h00000000000000000000000000000000, /* 3744 */
128'h00000000000000000000000000000000, /* 3745 */
128'h00000000000000000000000000000000, /* 3746 */
128'h00000000000000000000000000000000, /* 3747 */
128'h00000000000000000000000000000000, /* 3748 */
128'h00000000000000000000000000000000, /* 3749 */
128'h00000000000000000000000000000000, /* 3750 */
128'h00000000000000000000000000000000, /* 3751 */
128'h00000000000000000000000000000000, /* 3752 */
128'h00000000000000000000000000000000, /* 3753 */
128'h00000000000000000000000000000000, /* 3754 */
128'h00000000000000000000000000000000, /* 3755 */
128'h00000000000000000000000000000000, /* 3756 */
128'h00000000000000000000000000000000, /* 3757 */
128'h00000000000000000000000000000000, /* 3758 */
128'h00000000000000000000000000000000, /* 3759 */
128'h00000000000000000000000000000000, /* 3760 */
128'h00000000000000000000000000000000, /* 3761 */
128'h00000000000000000000000000000000, /* 3762 */
128'h00000000000000000000000000000000, /* 3763 */
128'h00000000000000000000000000000000, /* 3764 */
128'h00000000000000000000000000000000, /* 3765 */
128'h00000000000000000000000000000000, /* 3766 */
128'h00000000000000000000000000000000, /* 3767 */
128'h00000000000000000000000000000000, /* 3768 */
128'h00000000000000000000000000000000, /* 3769 */
128'h00000000000000000000000000000000, /* 3770 */
128'h00000000000000000000000000000000, /* 3771 */
128'h00000000000000000000000000000000, /* 3772 */
128'h00000000000000000000000000000000, /* 3773 */
128'h00000000000000000000000000000000, /* 3774 */
128'h00000000000000000000000000000000, /* 3775 */
128'h00000000000000000000000000000000, /* 3776 */
128'h00000000000000000000000000000000, /* 3777 */
128'h00000000000000000000000000000000, /* 3778 */
128'h00000000000000000000000000000000, /* 3779 */
128'h00000000000000000000000000000000, /* 3780 */
128'h00000000000000000000000000000000, /* 3781 */
128'h00000000000000000000000000000000, /* 3782 */
128'h00000000000000000000000000000000, /* 3783 */
128'h00000000000000000000000000000000, /* 3784 */
128'h00000000000000000000000000000000, /* 3785 */
128'h00000000000000000000000000000000, /* 3786 */
128'h00000000000000000000000000000000, /* 3787 */
128'h00000000000000000000000000000000, /* 3788 */
128'h00000000000000000000000000000000, /* 3789 */
128'h00000000000000000000000000000000, /* 3790 */
128'h00000000000000000000000000000000, /* 3791 */
128'h00000000000000000000000000000000, /* 3792 */
128'h00000000000000000000000000000000, /* 3793 */
128'h00000000000000000000000000000000, /* 3794 */
128'h00000000000000000000000000000000, /* 3795 */
128'h00000000000000000000000000000000, /* 3796 */
128'h00000000000000000000000000000000, /* 3797 */
128'h00000000000000000000000000000000, /* 3798 */
128'h00000000000000000000000000000000, /* 3799 */
128'h00000000000000000000000000000000, /* 3800 */
128'h00000000000000000000000000000000, /* 3801 */
128'h00000000000000000000000000000000, /* 3802 */
128'h00000000000000000000000000000000, /* 3803 */
128'h00000000000000000000000000000000, /* 3804 */
128'h00000000000000000000000000000000, /* 3805 */
128'h00000000000000000000000000000000, /* 3806 */
128'h00000000000000000000000000000000, /* 3807 */
128'h00000000000000000000000000000000, /* 3808 */
128'h00000000000000000000000000000000, /* 3809 */
128'h00000000000000000000000000000000, /* 3810 */
128'h00000000000000000000000000000000, /* 3811 */
128'h00000000000000000000000000000000, /* 3812 */
128'h00000000000000000000000000000000, /* 3813 */
128'h00000000000000000000000000000000, /* 3814 */
128'h00000000000000000000000000000000, /* 3815 */
128'h00000000000000000000000000000000, /* 3816 */
128'h00000000000000000000000000000000, /* 3817 */
128'h00000000000000000000000000000000, /* 3818 */
128'h00000000000000000000000000000000, /* 3819 */
128'h00000000000000000000000000000000, /* 3820 */
128'h00000000000000000000000000000000, /* 3821 */
128'h00000000000000000000000000000000, /* 3822 */
128'h00000000000000000000000000000000, /* 3823 */
128'h00000000000000000000000000000000, /* 3824 */
128'h00000000000000000000000000000000, /* 3825 */
128'h00000000000000000000000000000000, /* 3826 */
128'h00000000000000000000000000000000, /* 3827 */
128'h00000000000000000000000000000000, /* 3828 */
128'h00000000000000000000000000000000, /* 3829 */
128'h00000000000000000000000000000000, /* 3830 */
128'h00000000000000000000000000000000, /* 3831 */
128'h00000000000000000000000000000000, /* 3832 */
128'h00000000000000000000000000000000, /* 3833 */
128'h00000000000000000000000000000000, /* 3834 */
128'h00000000000000000000000000000000, /* 3835 */
128'h00000000000000000000000000000000, /* 3836 */
128'h00000000000000000000000000000000, /* 3837 */
128'h00000000000000000000000000000000, /* 3838 */
128'h00000000000000000000000000000000, /* 3839 */
128'h00000000000000000000000000000000, /* 3840 */
128'h00000000000000000000000000000000, /* 3841 */
128'h00000000000000000000000000000000, /* 3842 */
128'h00000000000000000000000000000000, /* 3843 */
128'h00000000000000000000000000000000, /* 3844 */
128'h00000000000000000000000000000000, /* 3845 */
128'h00000000000000000000000000000000, /* 3846 */
128'h00000000000000000000000000000000, /* 3847 */
128'h00000000000000000000000000000000, /* 3848 */
128'h00000000000000000000000000000000, /* 3849 */
128'h00000000000000000000000000000000, /* 3850 */
128'h00000000000000000000000000000000, /* 3851 */
128'h00000000000000000000000000000000, /* 3852 */
128'h00000000000000000000000000000000, /* 3853 */
128'h00000000000000000000000000000000, /* 3854 */
128'h00000000000000000000000000000000, /* 3855 */
128'h00000000000000000000000000000000, /* 3856 */
128'h00000000000000000000000000000000, /* 3857 */
128'h00000000000000000000000000000000, /* 3858 */
128'h00000000000000000000000000000000, /* 3859 */
128'h00000000000000000000000000000000, /* 3860 */
128'h00000000000000000000000000000000, /* 3861 */
128'h00000000000000000000000000000000, /* 3862 */
128'h00000000000000000000000000000000, /* 3863 */
128'h00000000000000000000000000000000, /* 3864 */
128'h00000000000000000000000000000000, /* 3865 */
128'h00000000000000000000000000000000, /* 3866 */
128'h00000000000000000000000000000000, /* 3867 */
128'h00000000000000000000000000000000, /* 3868 */
128'h00000000000000000000000000000000, /* 3869 */
128'h00000000000000000000000000000000, /* 3870 */
128'h00000000000000000000000000000000, /* 3871 */
128'h00000000000000000000000000000000, /* 3872 */
128'h00000000000000000000000000000000, /* 3873 */
128'h00000000000000000000000000000000, /* 3874 */
128'h00000000000000000000000000000000, /* 3875 */
128'h00000000000000000000000000000000, /* 3876 */
128'h00000000000000000000000000000000, /* 3877 */
128'h00000000000000000000000000000000, /* 3878 */
128'h00000000000000000000000000000000, /* 3879 */
128'h00000000000000000000000000000000, /* 3880 */
128'h00000000000000000000000000000000, /* 3881 */
128'h00000000000000000000000000000000, /* 3882 */
128'h00000000000000000000000000000000, /* 3883 */
128'h00000000000000000000000000000000, /* 3884 */
128'h00000000000000000000000000000000, /* 3885 */
128'h00000000000000000000000000000000, /* 3886 */
128'h00000000000000000000000000000000, /* 3887 */
128'h00000000000000000000000000000000, /* 3888 */
128'h00000000000000000000000000000000, /* 3889 */
128'h00000000000000000000000000000000, /* 3890 */
128'h00000000000000000000000000000000, /* 3891 */
128'h00000000000000000000000000000000, /* 3892 */
128'h00000000000000000000000000000000, /* 3893 */
128'h00000000000000000000000000000000, /* 3894 */
128'h00000000000000000000000000000000, /* 3895 */
128'h00000000000000000000000000000000, /* 3896 */
128'h00000000000000000000000000000000, /* 3897 */
128'h00000000000000000000000000000000, /* 3898 */
128'h00000000000000000000000000000000, /* 3899 */
128'h00000000000000000000000000000000, /* 3900 */
128'h00000000000000000000000000000000, /* 3901 */
128'h00000000000000000000000000000000, /* 3902 */
128'h00000000000000000000000000000000, /* 3903 */
128'h00000000000000000000000000000000, /* 3904 */
128'h00000000000000000000000000000000, /* 3905 */
128'h00000000000000000000000000000000, /* 3906 */
128'h00000000000000000000000000000000, /* 3907 */
128'h00000000000000000000000000000000, /* 3908 */
128'h00000000000000000000000000000000, /* 3909 */
128'h00000000000000000000000000000000, /* 3910 */
128'h00000000000000000000000000000000, /* 3911 */
128'h00000000000000000000000000000000, /* 3912 */
128'h00000000000000000000000000000000, /* 3913 */
128'h00000000000000000000000000000000, /* 3914 */
128'h00000000000000000000000000000000, /* 3915 */
128'h00000000000000000000000000000000, /* 3916 */
128'h00000000000000000000000000000000, /* 3917 */
128'h00000000000000000000000000000000, /* 3918 */
128'h00000000000000000000000000000000, /* 3919 */
128'h00000000000000000000000000000000, /* 3920 */
128'h00000000000000000000000000000000, /* 3921 */
128'h00000000000000000000000000000000, /* 3922 */
128'h00000000000000000000000000000000, /* 3923 */
128'h00000000000000000000000000000000, /* 3924 */
128'h00000000000000000000000000000000, /* 3925 */
128'h00000000000000000000000000000000, /* 3926 */
128'h00000000000000000000000000000000, /* 3927 */
128'h00000000000000000000000000000000, /* 3928 */
128'h00000000000000000000000000000000, /* 3929 */
128'h00000000000000000000000000000000, /* 3930 */
128'h00000000000000000000000000000000, /* 3931 */
128'h00000000000000000000000000000000, /* 3932 */
128'h00000000000000000000000000000000, /* 3933 */
128'h00000000000000000000000000000000, /* 3934 */
128'h00000000000000000000000000000000, /* 3935 */
128'h00000000000000000000000000000000, /* 3936 */
128'h00000000000000000000000000000000, /* 3937 */
128'h00000000000000000000000000000000, /* 3938 */
128'h00000000000000000000000000000000, /* 3939 */
128'h00000000000000000000000000000000, /* 3940 */
128'h00000000000000000000000000000000, /* 3941 */
128'h00000000000000000000000000000000, /* 3942 */
128'h00000000000000000000000000000000, /* 3943 */
128'h00000000000000000000000000000000, /* 3944 */
128'h00000000000000000000000000000000, /* 3945 */
128'h00000000000000000000000000000000, /* 3946 */
128'h00000000000000000000000000000000, /* 3947 */
128'h00000000000000000000000000000000, /* 3948 */
128'h00000000000000000000000000000000, /* 3949 */
128'h00000000000000000000000000000000, /* 3950 */
128'h00000000000000000000000000000000, /* 3951 */
128'h00000000000000000000000000000000, /* 3952 */
128'h00000000000000000000000000000000, /* 3953 */
128'h00000000000000000000000000000000, /* 3954 */
128'h00000000000000000000000000000000, /* 3955 */
128'h00000000000000000000000000000000, /* 3956 */
128'h00000000000000000000000000000000, /* 3957 */
128'h00000000000000000000000000000000, /* 3958 */
128'h00000000000000000000000000000000, /* 3959 */
128'h00000000000000000000000000000000, /* 3960 */
128'h00000000000000000000000000000000, /* 3961 */
128'h00000000000000000000000000000000, /* 3962 */
128'h00000000000000000000000000000000, /* 3963 */
128'h00000000000000000000000000000000, /* 3964 */
128'h00000000000000000000000000000000, /* 3965 */
128'h00000000000000000000000000000000, /* 3966 */
128'h00000000000000000000000000000000, /* 3967 */
128'h00000000000000000000000000000000, /* 3968 */
128'h00000000000000000000000000000000, /* 3969 */
128'h00000000000000000000000000000000, /* 3970 */
128'h00000000000000000000000000000000, /* 3971 */
128'h00000000000000000000000000000000, /* 3972 */
128'h00000000000000000000000000000000, /* 3973 */
128'h00000000000000000000000000000000, /* 3974 */
128'h00000000000000000000000000000000, /* 3975 */
128'h00000000000000000000000000000000, /* 3976 */
128'h00000000000000000000000000000000, /* 3977 */
128'h00000000000000000000000000000000, /* 3978 */
128'h00000000000000000000000000000000, /* 3979 */
128'h00000000000000000000000000000000, /* 3980 */
128'h00000000000000000000000000000000, /* 3981 */
128'h00000000000000000000000000000000, /* 3982 */
128'h00000000000000000000000000000000, /* 3983 */
128'h00000000000000000000000000000000, /* 3984 */
128'h00000000000000000000000000000000, /* 3985 */
128'h00000000000000000000000000000000, /* 3986 */
128'h00000000000000000000000000000000, /* 3987 */
128'h00000000000000000000000000000000, /* 3988 */
128'h00000000000000000000000000000000, /* 3989 */
128'h00000000000000000000000000000000, /* 3990 */
128'h00000000000000000000000000000000, /* 3991 */
128'h00000000000000000000000000000000, /* 3992 */
128'h00000000000000000000000000000000, /* 3993 */
128'h00000000000000000000000000000000, /* 3994 */
128'h00000000000000000000000000000000, /* 3995 */
128'h00000000000000000000000000000000, /* 3996 */
128'h00000000000000000000000000000000, /* 3997 */
128'h00000000000000000000000000000000, /* 3998 */
128'h00000000000000000000000000000000, /* 3999 */
128'h00000000000000000000000000000000, /* 4000 */
128'h00000000000000000000000000000000, /* 4001 */
128'h00000000000000000000000000000000, /* 4002 */
128'h00000000000000000000000000000000, /* 4003 */
128'h00000000000000000000000000000000, /* 4004 */
128'h00000000000000000000000000000000, /* 4005 */
128'h00000000000000000000000000000000, /* 4006 */
128'h00000000000000000000000000000000, /* 4007 */
128'h00000000000000000000000000000000, /* 4008 */
128'h00000000000000000000000000000000, /* 4009 */
128'h00000000000000000000000000000000, /* 4010 */
128'h00000000000000000000000000000000, /* 4011 */
128'h00000000000000000000000000000000, /* 4012 */
128'h00000000000000000000000000000000, /* 4013 */
128'h00000000000000000000000000000000, /* 4014 */
128'h00000000000000000000000000000000, /* 4015 */
128'h00000000000000000000000000000000, /* 4016 */
128'h00000000000000000000000000000000, /* 4017 */
128'h00000000000000000000000000000000, /* 4018 */
128'h00000000000000000000000000000000, /* 4019 */
128'h00000000000000000000000000000000, /* 4020 */
128'h00000000000000000000000000000000, /* 4021 */
128'h00000000000000000000000000000000, /* 4022 */
128'h00000000000000000000000000000000, /* 4023 */
128'h00000000000000000000000000000000, /* 4024 */
128'h00000000000000000000000000000000, /* 4025 */
128'h00000000000000000000000000000000, /* 4026 */
128'h00000000000000000000000000000000, /* 4027 */
128'h00000000000000000000000000000000, /* 4028 */
128'h00000000000000000000000000000000, /* 4029 */
128'h00000000000000000000000000000000, /* 4030 */
128'h00000000000000000000000000000000, /* 4031 */
128'h00000000000000000000000000000000, /* 4032 */
128'h00000000000000000000000000000000, /* 4033 */
128'h00000000000000000000000000000000, /* 4034 */
128'h00000000000000000000000000000000, /* 4035 */
128'h00000000000000000000000000000000, /* 4036 */
128'h00000000000000000000000000000000, /* 4037 */
128'h00000000000000000000000000000000, /* 4038 */
128'h00000000000000000000000000000000, /* 4039 */
128'h00000000000000000000000000000000, /* 4040 */
128'h00000000000000000000000000000000, /* 4041 */
128'h00000000000000000000000000000000, /* 4042 */
128'h00000000000000000000000000000000, /* 4043 */
128'h00000000000000000000000000000000, /* 4044 */
128'h00000000000000000000000000000000, /* 4045 */
128'h00000000000000000000000000000000, /* 4046 */
128'h00000000000000000000000000000000, /* 4047 */
128'h00000000000000000000000000000000, /* 4048 */
128'h00000000000000000000000000000000, /* 4049 */
128'h00000000000000000000000000000000, /* 4050 */
128'h00000000000000000000000000000000, /* 4051 */
128'h00000000000000000000000000000000, /* 4052 */
128'h00000000000000000000000000000000, /* 4053 */
128'h00000000000000000000000000000000, /* 4054 */
128'h00000000000000000000000000000000, /* 4055 */
128'h00000000000000000000000000000000, /* 4056 */
128'h00000000000000000000000000000000, /* 4057 */
128'h00000000000000000000000000000000, /* 4058 */
128'h00000000000000000000000000000000, /* 4059 */
128'h00000000000000000000000000000000, /* 4060 */
128'h00000000000000000000000000000000, /* 4061 */
128'h00000000000000000000000000000000, /* 4062 */
128'h00000000000000000000000000000000, /* 4063 */
128'h00000000000000000000000000000000, /* 4064 */
128'h00000000000000000000000000000000, /* 4065 */
128'h00000000000000000000000000000000, /* 4066 */
128'h00000000000000000000000000000000, /* 4067 */
128'h00000000000000000000000000000000, /* 4068 */
128'h00000000000000000000000000000000, /* 4069 */
128'h00000000000000000000000000000000, /* 4070 */
128'h00000000000000000000000000000000, /* 4071 */
128'h00000000000000000000000000000000, /* 4072 */
128'h00000000000000000000000000000000, /* 4073 */
128'h00000000000000000000000000000000, /* 4074 */
128'h00000000000000000000000000000000, /* 4075 */
128'h00000000000000000000000000000000, /* 4076 */
128'h00000000000000000000000000000000, /* 4077 */
128'h00000000000000000000000000000000, /* 4078 */
128'h00000000000000000000000000000000, /* 4079 */
128'h00000000000000000000000000000000, /* 4080 */
128'h00000000000000000000000000000000, /* 4081 */
128'h00000000000000000000000000000000, /* 4082 */
128'h00000000000000000000000000000000, /* 4083 */
128'h00000000000000000000000000000000, /* 4084 */
128'h00000000000000000000000000000000, /* 4085 */
128'h00000000000000000000000000000000, /* 4086 */
128'h00000000000000000000000000000000, /* 4087 */
128'h00000000000000000000000000000000, /* 4088 */
128'h00000000000000000000000000000000, /* 4089 */
128'h00000000000000000000000000000000, /* 4090 */
128'h00000000000000000000000000000000, /* 4091 */
128'h00000000000000000000000000000000, /* 4092 */
128'h00000000000000000000000000000000, /* 4093 */
128'h00000000000000000000000000000000, /* 4094 */
128'h00000000000000000000000000000000  /* 4095 */
    };

   logic [BRAM_ADDR_BLK_BITS-1:0] ram_block_addr, ram_block_addr_delay;
   logic [BRAM_ADDR_LSB_BITS-1:0] ram_lsb_addr, ram_lsb_addr_delay;
   logic [BRAM_WIDTH/8-1:0]       ram_we_full;
   logic [BRAM_WIDTH-1:0]         ram_wrdata_full, ram_rddata_full;
   int                            ram_rddata_shift, ram_we_shift;

   assign ram_block_addr = addr_i >> BRAM_ADDR_LSB_BITS + BRAM_OFFSET_BITS;
   assign ram_lsb_addr = addr_i >> BRAM_OFFSET_BITS;
   assign ram_we_shift = ram_lsb_addr << BRAM_OFFSET_BITS; // avoid ISim error
   assign ram_we_full = ram_we << ram_we_shift;
   assign ram_wrdata_full = {(BRAM_WIDTH / 64){wdata_i}};

   always @(posedge clk_i)
    begin
     if (req_i) begin
        ram_block_addr_delay <= ram_block_addr;
        ram_lsb_addr_delay <= ram_lsb_addr;
        foreach (ram_we_full[i])
          if(ram_we_full[i]) ram[ram_block_addr][i*8 +:8] <= ram_wrdata_full[i*8 +: 8];
     end
    end

   assign ram_rddata_full = ram[ram_block_addr_delay];
   assign ram_rddata_shift = ram_lsb_addr_delay << (BRAM_OFFSET_BITS + 3); // avoid ISim error
   assign rdata_o = ram_rddata_full >> ram_rddata_shift;

endmodule


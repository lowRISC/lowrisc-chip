`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jV86F9yDZRipVbWW+/Be9dUIvO1203e0/QSaJAwx2llqLHjiQPFnp4sI2fcmymvV7wbHazAkDZgw
JS7+xOzSR18VfM1G7uj9WA4HA2f4t7Rf5q5Uwg6AuRgGRcdKhzqTuyy6XSJ5jn299H19qQxTHlMB
xs4CmDV06QXz+N1us2mVCuPG56srvhqcqnxXNOqXvvvoP67BLGfO0Gm+7w1/tSA7WVrCRZO6f+EU
H0+AXuAOOrj7LRqPDZn2zYtPALJH6A1HRioZy7HoLRpJgRlVzCGz21czZnxTmeF2jC7iWn3UQVG4
4/LGuca8S1huB4TZDclR21PKUWIGXr4boS8/dQ==

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
PDB5hU5vy7YI/dpXUPo99a/WaBcWlwFeziOAK5DiRaioIQrdo9xiQ4TXkP17N1rufAjEuxvYpC9b
Wyzf7WvKyQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TMhFzfm/qsk/dJ3AX0Z/JaHeIz5WOuqqOuRuF+TrajePXy9T7MOAiZG0858t6BLImZ7KF9JAZUdb
sHhmy81vatWvE9Ig7nT3xsW8Sg/eJQotm3jdGDbBSK6An7AR8kLagTrt7aSG6bAn8lcQv4ciBwfj
3yaMsw5ZiMJLX/y7NaI=

`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aIZiJXiyjnjWO+9L9VFEo7qsa7a8wtRX7khE7jIaXquFxJ/68AOQ8YPR64aoYdhHjWpWGYr82fgo
1O6ucjko82cPgKb4larmI0uh4ZVfmtAIPwKrIzA5nqHeNjlMrDYf7x9efYLzwkGTUtuedDlgblc8
RFQjObyh5GCv03NolVM=

`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YRFu3VWNK/y4aqaWwxub+hggoscun+8Oo4Z7PgLf1jcrVBr3TyQivMFnWGEcMmdK5eKurw6sgRqm
X5xM6tNTM1xbRMoqj32DpB1/luNKjXMlwT5mKH8wTz9Izk2Qr/2rPsm8wtJZ6o6NIHDcYa4+gyG9
yEYnlDlhEOc34+r5y/DpoKQrZai3Ku+PUFV5pAfFWGRozP5TAPLF3PQ2ZsE9XIvg50XAG7f0DNhJ
VoGMYAIIaw9Uw1QL6Iy11XdvywXAZG+Uhr+OxlfagmqpF3SujK1hwDc/hEARQPGoXcs2t7kYsCgi
qhABkl3NVrF3AC6YrN8CowfR5AHUmjyaRfULqA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15024)
`pragma protect data_block
rWrlwpnLj89zhtcaP82+sdYPWqNoFGFOKl30QenCr08EBVjzDuiyeNNqsJV6qszGPwKdrd1M+ID7
UERS5MkRu6Fe/eBipWhmWu0wybvnw1/YDpd32ZB/rU/PrIC8QUf1Zoxpwk2RBBZDEmmRxWDBz0Pn
0oN5nHe5bRCHjUzw937aQIhtQtUjrpTshpkmKaqGsZI6Uwzp6GCD2v/yGZ/+8Fd1NkgP0FClYN+y
igEPyS1W5HFWAlj4MXpwfB0TtftO7weHFH+QF+9nql4BDcCZ/5dPaAGLL/hwf8PzCbjXbkfk8UQz
h8Z6seSKhRrz+LxKRUdgKsekoOr9Lyj4Hff2kiU6/U4ZrzE/MOm+MAyCNgZagegFSdM88iDQh/8n
vL+OcZ7Vi5+YN/NCoDEaW+NndBL5FRbVs/37/nUH1371KHAmxxQDckKjvCCpSl2FuEwNWq7ESggs
X8TjPmN0gmbHBOa12mrOpjgq5iDhh/Va7SqkYg2uVTA+lp3gVbI5vS0UGb6kJAMgL+oMeV8MVktP
ayi+p0BYHlLfqiTUldkTxCqwCGQPw3vf5AIKvX3ZRy0FEkGJq0bnWlKsUZjpq8zvXKxgCm5in3zK
AqAVK6Dsenu/ekyogpKogunwWSBW8ELeuwOVbSadzYzVf2X1FmUh7/lBv80ZWhwER3nmLRbIgPVH
jxsegl/YAAkVlVShL+nqYxIqin1Gfyxe9So2MGw9kAWuX0g/732+pCH4J7UPpYHJPn9onFsgSqQZ
x96xXaDJiNglZjUk2jOyTUqqFSpaBINYhcOc2x1F8BLcDv74AnHAzcSrNu0O2bnBO843Msc9EDRP
LOR8PhWrXFkfHzq9egv+cUgmg9h7IYzZu8dBkkfKtuGvjyFXNxYIPWQD17es5T+8N7Nx6pWE/my8
pZVILmFj32VKF4zLusjCcSF5cnALFMw7q64G62QFHbc1l9eh0A6VtYtMqM9c4Cg9wQhnCzQszR5P
ekgfUuuVVv4cyej387B2PFY/591TBWvSYuzP4MCNSVOgJjuME9XwzluUgMuL51X5oSedWCXw6z6U
0aoB0gVG2Siqg/K2p5qNgaZNmk8SAGgPcGOohPFFiWlzGnwhFTYwDLmXhrCIDK8vUPkdYJrG8W3Z
yX55ARig7aVpOwHtAny//r56IeefpZTIa9wT+lbUJ6AR2wRThIdYlXVOz8N0quAoMq9hRRowq37+
F+CxoP155Bjo7/XBpsuB0KbnFFdkiFw1Jl1+TwwFHcVWpu2BvxzPYZXeJ0UUZD4P+g8ndwgK3a2a
t3zD10ZmlZl44Lsd8ust9Hw3QmDJMHX7ZExZDXVCHMyeRWXQWFskwWY0LqlmFx+XqSQcMc6emD3H
grb2e8VCRsWaDbRQG2vcC3W1H8ba2n5zDG62V+ULMbkoTxB+YyRSn8R5dQ+nEyPI0jsAAYpDFP8A
IowOfNnZNEqGcBv4ebzFs/ODoxs1MtWjCk0Qoeh3retIsVrCFCAIlN2qZazj9PGcE3kSzGcjQnMb
qMUjh8q+G0X8AB2pSu9ezglzAfbbj+QfYaosC5mJ9WKwVCOqFh9UHaTYnuJSg2mKoNxAxV41Hz56
aQiWRlOgtZjahV0dPo1KTilxJOLrn3prFFsE7AcJQFjLgMU5h2venVak0VUpIr3N0UidiQ3Ocoor
7ovxMKjqI1QhGzcFfWkU+ynJqeLziBeysMOmfJtWLvPuZeESu0i38LERj6SCY7eu3W5k/3rB2rNg
lidYOA5tfXh0UdG8VPN/TjU9GIVm5x1pUdb8qPywPiupO037B2OjxvQ+y6IGd8AXBXGo3d1qM/mn
uQz1CGY4PNBAkn3vEn7PR2b9bqCK0BaEgP4MQUWtPe0JdZxnf+6tuex9bJrf46dBxpfHOoOWfHVy
AhSevLFtVuUp1bBnpmOfjDIYJyyAuUQ/kofq3xnVnYVKs1Ntwe+nBmNu1qm+GbRjJXq1SPNHcNhD
8zB9mKI5qTD7twvPZ2ZsRsb364ikFqRDM/Mw99kbdzL7Q7vnKHRf6yDaxlhXu8Aw5VLJ4gtpq4yL
VJpvN1bLShaYLmS4R7995j69yitkUQxww0pAzUcfQJTUlK/CE3R1rRrwh7sDQtYxB2Uqua0WE8fN
507EOIG09QDlpV69qUSDmSHzTSIYhoDV7tAHIwVQPS/ro+4OCWOnBAkj2+VgwuQ/3q0NwX88kiOc
9HbgXotI+NXO6GSjnCJXEVb2VCR3OwQKeF/809+iM9BMx6a1youkDiCwHn9rqkSAVvlS6OSiJllh
WkRgll+9g1kxSXSdQsYtzeryDZSNlqt3jGr4WPcSyDoUA0LSYWY2y2/EcMPCTbpoCWia9giu4INs
KAol9/fkRtwyRFSLKkEP6ubJJsOnzC6D476m9++ripHQRxQcgGTlvokc9nhpTCq1jFbprxk6i0aV
fx+WdLoTo2KjrzyWoWyJ132+9FdJ26M8kOWkGvZHoyxh8bn4RWUHSwkfkDrLeCW3sax3ND90rxYY
Xxsh7+7rZIktFt/1bM/AAF0KYJVv/g+xxR8qX9vBN/fGT6H4aZn4Dx8wTSA8nYSfxtd3L4FZt1dZ
Uqa5CHlS81Qmrbv3sw2J8UydXTwqEGsivjiqlwcyb/wHMi5vZdhnfSjmXCcgvcaLqoR+lDPkjYrQ
5XZbZl7iqGCGwMccRztvTz0oYOF182voHqqwcw+9Poun3XMW971942n/P1j8HRaAaKVrPOJRiz1K
BEg8P1wu9UcZyIsdlzIBlTkd0Hl38InAvyf4dXcHbigkPq9/lYctOdIV52KROdC+0e5mTgUN9ZQX
KMLyvjgmKQMijbninnxSAGWHqAMfUtyzylOTfii2vPdcAZbFDDkKolWGv64APpluoTfvTtuVbLO9
itU84X0DTRhml70bnbK0qHHLHig7r930Hg1IR1/Y6KgWuiFqT+7LgERjzjoo2e7wXcq8Hz/yF4dR
p2ZLgVkMSLYlpFjBUn4dn7OrvzIXV8cijIMvokYL0LF7UbUlT4SIi0+i2Vf52U14PUw+pISLnD6Y
l9DhNUvH6IKWjhCPG/HJTyyKCcgcAjNFBGREXJwuVZVI2bl7AgWnHhKWSkaDnCy3/QV2CKdmzatC
UC+8hXpSFDPhgoL10JrPqrWrYHx2gTwi1M/KQrBmZ/CUopGWiq9f7Kzu6wgEnwP3K3ySQQo3jSm5
b2Y4zVq25p2/5lEsw6fa6pZ6XAKunplcVao5tU+k7LO1LMnOM4EmL3sb7dsZ7hOenzJQN4+zCC/j
aoHjzK9FRjz1TMUmJuO8ahP72tk3saQQYPsXThqWbc+8F4uorGpywwVsMCKQbZg6lJzzoP+ctNcs
Z/4TqdbNSXrqFcXuVv6eljzZrxbYMVpRFeaD27JZ+YrtZUcIzI/qhIjCbhfzJHvCPuQXW4NRwqpb
G2pbrcDrswoIWQzgoyWwRs5WifjvOOLmMvBTPz/7r5O92mTJTKhM7wEoEP9ZbnDfsIHfpTHbIslz
Be2bPpuLR8HPleFgi1XJn1xsnFVXb2uBvSdZvu1JAw00TvQWO92KM+0j5Yohmbi4809htmx8C9yy
zDAB4PLujTaaKzJXCwiFzQZ4R8IVTSUkOlce+Rl+5S4xBRw4/FM1c1Y2GlGjfouOmvjGY56vg5+/
5tBEk8+c7HILzL129LAd8v7qMBhXHz12wZy9nipthgfPJHirIxY4wTKKxhfc6/dnyS7N+K/hUrbB
iMpXjKY67rrJxMcHL8d9cawmW7YDoK5UqVVPXDG81hGhtlnN3Ydatm22Q2bTs05TcR0TuODVXXaY
CDVYCPlV9G/duyhUPpliEO3GhBuXr8/5cbAdSyQcNxBp7cFvWjWPS9gdZoc18YbLO/MkmmsiJuse
qPH9XswvHmiEe+WtbICFqNlIiNwboTybtK/nUvu6EEdIJnijH4wPEAgtzKVQuiZvXcZylwus7SDZ
vv6h6HJuaAynpWaZIwbTRk6aBQVyPQYN04YSAIvUroyfPgbJwePJhVOR78kXSSPY1FCvcB3MS9r3
jI16iB0fvanHSmjGNVQ3xDyyJXKUUyI88UmllgrUuTZtj9pHFKnJIBUt0FmFtCqJ1VDQFfgxstzD
6uuIC72GRPgiltpuG2MFQ9LzpmiPzR2TCzKQF79w7X1fyQZHjztaQgzW32WpPnoNyZNbfCRmozXl
R8lA+KcJFKGRYZNJm5NVlBY+eJSrQvh5gcEPlN7UrbL9cFBDIGYX6wHbSYQzS+vptmUjxt+Ff8nI
X/NYWdPMdsTaVstjEgthuHSZrzs8Lj0mqKotdPyROczuTMIXTm+EyBnQTFfdOcEIZlQ3BTeppb5O
N0yuyQgOzl98iWYsc7z0pVKe2xRkR8VPd7Ii2porMwazazuZQb/4sOQil7C9TAbAJb1ChebTZcA8
IYIxR0d9bcV8itwkIrPw9m5GEVoCEI2Kw6vihFr+/+lfAtlResUUqXh0EMHLnJxno2fVh/mFnErx
OrzmSJmN+XygMyODGpMac07fTOE62QgijsKO6LpFDvUIpNhCOGbJZfc29knCRiVvq7oTV8RIvrHg
ZNDEj1H6/KAYkRxIfNfIdRNEGM43na1UkEjUP3reoL0IoaD5tG5/AFeWUixuDinnztuMgVksyWoY
cgSvUFkSrkEubnR2OT+BH/fdDJB9+1RrBKXlVo5ZxMM4Y9ZDxhEf0qX4+LhYZsQnUDlXoVBCvbNH
dlQFVqnPMSQCUMQ2Ms8hQgzkKJWdPJoJnp71gEYuAnQ+shtvu1YEd9ynYR+HnTNjMK837zAhG7uM
bmV6R8led22QBjk/NDi8WVi03+T5lmRKa9/ubLZbUiiY+5oNSIprZNfILSZKUVG2KMtVrgV43n5a
2ogMLaSwSmzgr+Deow70Pmt0AYZtVFsSJRI+MB00qDjavRQX4cN2KJMYE3y4RNohosWURXWfkY19
pq4wOmANabrJrV4W74R1K1Q0/w/oqHHiJvnn6jhLyQUGSxMHfkwjcfuaVA3z1Uzi1kBfMi1w5P6X
Vi88E96RKt2zj4AKZ2locE6utxni+3D4HBNf4yIwFRogKFPblP5BC78Qb5adn9Kuu7UinWrKwHF8
YBTg9tIuZ+vgDayKdTI1PYu9Xtjh7HKZQPiaULgEpfiTasLlEQcmitxakZ5nV2HUdBezRjYmvn9X
iAZP/sibsYiMKS2NuniZ5OLiNAiyHR7Hjc0MDMSlrABnS2kQM3jjJp2uFWuh+3j81sdOj4aeXEm6
4lA0kf+0WjeNEAc8HTh+kl8kPlejMBu/SP2dE+SvsKbjr7EbipIeD5HhSD8EfIvPM1VbLJVtZQOd
C24cgy7LIXK0XgsTz6Ovrx3Cl+6QigX2VhD7mo0ln0MxsRw7J8ppLX8sk/H9G967MwbQYQU0c448
drD4GDHKiezOK1DjISoTxYixBfqGP+KwVvz7B7f+dQjBRtoLh324o6iEEw4bwheIgUZpSwHmcFtv
wr5e9PkmdRqm7b+5Xsl+gcnE0zMs6oauaoyjKL1twML6gM1MFVjuxEAyhCHCN8u1GxSHsCcYbmtz
fE/zxPMew20gPxaT2VTqCjJBEDE0YnemqawdUsy//dDtDDK0GjPRUdpgBuNzQxHRR7uM3MW13HS5
HWfok65CH8gCAYemV4amRvto6SpzD6qvv+6WrzuEPUnqeVnOZP5uJxm3JfwDL1vCKrxGy6oygzB+
3u4Ev6/KpFDJ2HZduNesvQLyflLAmihbBB+AWnn/0zLs+L/1pX2qerJePOpm0VL0AGDF/F8TyWjG
ar7NoX09Qhe3B9ZNXWrh0nYxWWmHGHDMHDsRl9v6/174LRHU4zRVvUh4Qnuh+2u7HxxaJFXFvDYU
NAuyqvdPts10Njut4cmGv6p+MPwbW11y0huBb0q85yBJVE3TunmjVGkR29js8pNZu4mkI1mhIXK0
PW8NDrOABco1YF9GMFNhdN/tjn8RKOeEjpHJoOyKDB4lxomtIuxWVCXPOutSSwKCNKJmHw1g+S8Z
2irzv72uk6RkN4KmIFBe/vJH5E7oTeh88oMvfKVSPWPRk1WUysaMVqjhlBzL6rULQAF9FFotD0TH
r5tsIdVxCYQDiU/iQLaiah0TrfOdamq/ZLkJzeWCO0JRwAdCSCWS8DtM6lHaK4BeXyGo8b1+9kzV
2gRJbXXC73+g5c7qY0+z+8LWEdgqVQ0XKQb8OuE5wWrJuL2eSjDB5I6d5L5DxETNmXNBBsrmRoEe
OuHmUEtA6OPxCGBRE2APk0Pf5s2rGK0hAZVKwEdZARYGS4Lr54LaYUWGOyPoq5+BCPSBhUXayWFp
D/BLoidBKetKkSA0VfoYdN7iZKJGB/HdFN+yzh3EPb1Vgzn945guMopDGm7CWTwULl0lkUknjm7/
jy3jS91O9rLN16nNDpc89XpjbmttbPAog8toZ/fK5VBUzZuQQMzVTS55QMcBOAILIRScXtninohk
smvc++tziAr1LaI04dSTUJ3dOf4kpgCQ+86irNmR5wC9XJBoaUnDtXMrbTp1r4bSZNPYvZuw94RP
r4B7Y8ZRoSvH5hDP4CgTs16oqx+4ruER8ZdGrCqdb7Cdtbdac6rM/3PSorBPvn/23UV/V1p3/gTz
lqpSKeVa1hKY93FdMHw+AMxTYK3n8Q0ALgmrI2xcdb2dFNJ+PCbP61Q5Xcn6YenCaq0m3rwFw5SR
9oeEyg+GdmnGhEn36zZe1VFkp2gXK2xhpdXcfgOvR83roK8+ujca9DyefKqGfaogwgquxG6rlokW
Hwmo907B+j7pxVbx/xkdYK0qT9tXqyuztHhV1b7jWBmmPG43Uh2YfJr+aDAXHz4lTCxQiZkTmbiO
wEJuF9+0WyQiojub9yau0XVj5vYQrqXm3ciMaKFYxYCJSQ7/RXHWomEsGkrBAjfsWKxME1enHX7a
ywn3OvUMkbuK/1hPD9Izn5GzgTehNp/Woe3JJMdTwtC7+OtVmlkO+xcNrNYuQ1Da8nd0vDK2f49v
DvzggHbyiLupmC1sXgUOydEFf3KdwR/6VlR+P5jMDkPxrF6fwDzVbjwx+37kpTeK8z2R3v9h6nCq
VUPzlcGcZds2/8Q9QBOIHIUIB9p2CuZGxsu3rLYtANkcKusVe/oLwacvQpESndB6IpBoYRKn5p9p
EgSMiTelCoBLLPPxXkYHFxdP+v5mAcAPrgbLJX8iTX6oB77BdggPPs1Usx5fNRowFGpv4X+UtIb6
xN1Br3R5+fJbWN28L3VNSERBuNdMEqwfQxIqfvI+i8UWbY8ca9Grti0o6nJYOJ939tvR9YtB4Cas
68zTBVW9PkTJ+fDAeliAXjc3W8Pb9rt5CCu+ccT4O+kc8jfWhMo6mc7C7MHOY9m6ZvkTVZjKXk4y
xbukyk0SW2CnbB6QxlAl279GwiRSglTh7qCqGep2D2PNHMl++K26ScHg5AB3bPJEzxKSB97ff9fG
ZtHA9pqVtkye2Rg1Eg46q4OYdE3dOB7HulmyXNw7k9H+NTTfRExO7SbcGHmlrTaRVM3UVWUqRc1a
iIPt/Ds+coQWyrU9KIV+fm7PYSA75iv2YjGwMmPeiHAydI8UCaSj28GkaH9SWiraHSiAJOY0YWjw
2imB0vStYUJYsD4aR77sTRWquhteU84dSWWywT8lQC4B62mf+6/bhbzo619RtKRS+RrUbxRAWvG6
BX02FnydiuzNwgL+bD55sVSVrVkkAnmL446Gs8CO45y6R+5VxXgA6tYEVVg3Kawgh4JSj7NKok1Z
fJpx0DT3jwO84T/+zB07/AiWY15rN9oNhFb9lxNO2q9KiQu+Q9mxmExE98+P/uGeSPoiZFik9QDF
8AeAVBXqxtew0sdnN65MEUTyB83MWbjZkMmNX89Ktmg1hhuWbvzbrY+Ar5mHx4wsAyPmaAxbEG6q
qf301HxSRSZz5kIRZLJD9d8H6hxkcC9hOR8wzW9SQ9nGMweG9pg0fiV6IFw2gmDIi797uFLSAzAU
yLsgxX0/MVDi/AF+MHk2UrmOmRnexAIlKB/Ebnl/Rmv+1/9J0FqKDR7CSBdNyJaWboCWuajGK0jF
im95m3zh+nZqBmUz3AF98WlfjBWsSaTULFz34sPBWj/TRMciXBaw/2wwAWSGdxpZ6RpNStSGNTVo
fYN7WoMjcxnQrvrWn2H6IM98iTpw22exK2TMPP5X7ulpheC71piiO9/RDTg8eK6G4dSdKGf5qffX
hf8mellw0jI+63FpvWGT8o4WopvsVDo9eXkqFr0yW+Wdzzd0rGpdAI9Iwkjld24GhZcop4SaIgGt
1sTz5Ls04hcIOrYyDKqSFXwAzmBlHAor3c6uZDIY7gFv4mN7szrv7uOQ9ipBrjBEsf7BsVaCHOkN
4kLDXWZVL9b7kY41S58raORS18qU6rS5FuX7eHb9BLJjJii0YmH6d+d4Rxa30oKHk4bA2hunWg8y
oWnmCDjn6YwBchLZYONg/n1tY2WDRi2mql0RXGqZ7bzPukJX51xR2eEEDh/Zeqju1yoNYFjQrkMM
XOvl7iZJm3AQY+5+n5gwJKvSVPJMgGbpHJG4iDHNE/SIiOJKuMeMJcDZLeOUoanOUnUKSOQ4eywA
01T6kQAk7o0WJ8swRxYVqUMXAzDZTz6xPBUdGxWOwyPTZdQo10JguHTy6nSxmVJBNTmHProjar2W
7qDroMPMqQwtQFcytzmDX7vOStyqD10A2aAG7uwxVeqFZPkMZisRAI/vcXCm3mF0Jw42WJLH+a2t
svadUnT6r4h6M3283RYjm4BNS3F9YZd3McBvatdibPuyafjEZa940xkbBV+01ERg0SfIZ68NzTDL
eMXGdXFTrfxuA0SOxl6sO2dG6nZjx3kW/Vy0R1M/DUQfxe6MECGbxs3x4wMrNd8zVdlpkozcib6a
rq/y9uUkQyIfBe0omBi6kIjUVPC2HLGS7Derd+ytxH821+sA2e3TdUfVFH9xTYAL9etCsMsqXs3U
Ku1jVbKjHV5QHlMwktqZOiClmKfVFhPBBHsAzZ2sZ72ZtpzrK02MKhFiz9R+TKbE26HCWrMcjTZi
QSl3fPfP2nn1pY3kUYmTfJZaxmg+oNyl+dQOsRgkTz+/2b97Ndzu2N2DzHiZZoPz3AIW22+8u6VP
gtnphXoGsAmz64ajTmtMCbDUOjnC+pdDMjaSAHSc6EpecoJ7mGQCJX7CLMOvCx57mW4yXZ7W86im
EEOFy6rhY5Gf01XW+Cliq+o8iewc8ULnUodcnWZyj0t5bYqU/eE1etDzEbgrvJKJIJJu052DVsz1
HramxLBVv82+MjosdQRYT0BFxwAoC99m9VIe342VNu1z0OvbRcUnGxVubnEz9poNgp57cqWgfAuG
N8Hr5hP3SpnmAK4dwLEBnvAOvb1QCUFDqnkkjN4mGDqG1BZXOIEiIOuhYhvlftFNxQRVDGyTi3gI
uH6ZUnUrS0d1asjsT26rU+CpoOzN8PF+LdD9Yjzk/idNjoEdgWv1rOjjYtC6/QXOT14xYKhH5lNH
WgvuRZXHz/U7LU4JNTbvACPaQroSrOZEK1gTaTCXSfbhOWmpTz3qmzGdD9nnc4c6W6j8oW/P8U+H
dNsAfZVwtTOHSpyUN8oBwrWPq5zBEFMrtW60l2FAd0qtP6ANkeGR0c+QgOUxnfM+doCjrczF83Ym
r4KLak2Bmz2ZQIiB5/YpBT4NnMJzattNnerorZWTE2QbSkQURBPMv+mhLUxuO8S72tnNR6EnVkW6
jdJz+6foQ0ollSl4xhLnZPAPskjRyjcnXpjpp0mURVkTlDyd7yT2WO4+hUgjhtF0k/03aXFnxMC5
RtkZP9HX6iTxZgPAhqj0l/LrexrS/c24taDGibMhZig9dEqp3v9Bb99tv04efYbpwLIYQd+dJyqI
XFIo+48Y1JPcDC/8TFLT4akooZIfZim6X0cmQCp7y05LEnjYEOdc7wa4BgNwYPht/+WlCPTp47WV
+B84nPJ2lbj/tcxjjSG1vXd744eUDCSirpQxN15OL/ugPNy2E1yvRCv20pxH0AO8zZhxrFa3uXtI
ebQ/b8GaZ0RyrcjeN30zaGiCWkAeUN6CbjJ1KDqQGSX66Qg+zDIi9YKJkLeJmvSu9L6bziMt1uTp
zm90NQDQH7dP695r4748aUsz/cFqpLB94urCuUq+jCk+5EH/16epFw5uGgh31C4FAw5Mdu9OIepJ
bfBFaze+szia0Q1P2HMUAVS2R+nve8+mY96rekJ38z03d225F0YmGm9DRjVvk5iXUm10G7U+Nq21
LeIjr/aZY951Y91K1grOOsS3M376eCEpLn1b7WFw6UHLeTjI8feceeUzGC8sM5EDZ1iGzULyaQ6+
TtbKXqMkmVg5ny03aPP3lXdcMBN/lban23Zw8FxYglYjt7nALs/SeiiR/il2X42BGIOoNdpcQYwt
Hmhbph2odEh/61ee4lFpiLVf992IRy7d8031V5482Tfd5ZsE0XVQSeEeJ0B4Btogrf6ZGRk7Smy8
9I4grRuYe3PoMvd/QzjjbSAWvs2oWdZtFXz8W5an2dgJx2pd18CLoMAINY2zDKe0NnJpccCctoJu
x1GZAdJZkfVMmAEqxVd5+kYndfjZCyBw+WlYv7D0/pvK4SBad3tMbubpY7NupSsxT22H+iwPCcyQ
JlYY+GCbBwJfW/Sy7XYXV7Iyj/fe0aAtT22KF5utTwj9dyeFzDSGZGfjD++UPGKaqBQh3eufk9w4
wOgFPkgBjcdxxha2QtZr/pEndh2f+zAzCVQREbgBPZIc2u8rlxeyDExu3Itf0vb0n0UD0/MQT1wA
1Fsqk9mJ1MrNEV/0huS2fUif9ZLjY/2M4ar3XdtO89olF4R0hbNkQJtIoHCLVH49KpWrales5mrU
fNgxzMffctRIgJdN/qS1BFTo8W20DKMUAWIuJ0Fx0GtWPZL6O6Hn+ZxvKr98l8dS6dkjXTkDfOKB
9vNLj831co9rGMvHm+ZS4joQcDEY9VuDfKODBsK/iKPnxso3r3Qzj+ynRl+76QlzFPibpE6koAnN
3IXUwwIolAz4655K3m40NYbR7TwIXC41fZT7ZJxHr8aUgbWyZrx8nvweeoYD05C8k/XACAIoMXd1
IOwiuUFFDBPDKohgrkn1whVlkcz9sAU2gqYr1+rQ7zd/tGThOp9nsrkhYXrsi67cMyq0SRW83s8t
vclALtG5P7Brekd2wWz6HzXtlwBkoOJGF3hzzYXeJauhd9r306FZMS4mMcYQiPLv4sFkB9EHhM4/
lgiO8pPw+LGeiWCI/xV5emXdJoCdcip2Cm28+lIZIU6BsIfDQSDxTyewASCSR7WLaOuFlFonV+h8
Cgw92MpHbXnZTBMRBN6G2DVYQt582SDlvpxUZbCrG2j1Rr1nneuimaBsjKgmg3OgolWTSfoNN53s
E4dwgC0X0bIKeyuhR6APWP3XOzGYY8F2Y8f03PnsD0VhbM1UGFs5rtCTvODL1qbGkfXFovMZiz7y
eTbfWxtWbZt5BTt6rJS2LzKaIN9M3RNjRKZFdGGjo18N04fTh2e9BFepsAe36z2xNiCAOQGJ5Y4g
PWvQ0GOgBqXqLRFbajHrC9Uqq1KQ6DSxG5NUgW+FgDeCo0nO4xMDGhJa7i6L1cwckGYGzjkQdKtT
npbUGqivzh5SOvudVDvOcLEpmD5SzmKEtA4MoMq9D3EOHoNh31kD9oAxXxmwyVrZ/jbRscWtz1KV
xaAda3CV+0uGhMqBQL+ojVbxraD3/U7bbFYqt7SZJ16xDRLRH8zjYpQ6BxXxTQqs0J6n+yMFV/IU
geaq1+fEZWi3jO1OX85WUBRiMy5KnKlSU7jskaJJ0W6SrWJrnxd4nWoJGr2qN7s2jodkP29KsYuo
TC/pp0CtY8Tfy/VdjRm3RrB1Y3Xc7WIVZxgOqsv8UB8G4Ika1Xv6G6ge3NMz58US+g6FRlwdm3zf
3V1PsU60YNN5uzE5fZuHFAQU6JsqmYMDlUp4VFpGH79xX8YXGYD9q5IFGD7iYlCbz4tq4v6kAz9F
ymF9vRat8BDzXQBthmDCYWoXjyaRZdlMBwr7I02orS2ijZD7TBw/oIRXcdnfKxF1j8zYH70HpgkC
FML9wdJ+MKIqHc5JNt0PloiRs9hXQ1UGBKpoZXnIfH6FXQs6unFp4e/hU2jJnivJlRvKIqD6m3p0
VP/frBLKV+fAIRpKNEKlUF6vPmMYJ3PXxQ4d+iGq9Q5WR3c6wx75USyOJloCrGywfYzd/nhRzbQv
uF7al0fiFlomTw3rZsVnCGwVR/RlaUErM6zkuRLAQ6/PEaB6P7mOwGZzUjX/DYkDeqdTr17+2gDm
tkbAR0g/0EdP+hsDwtAEOAFEBUeRe2BlwEIKmnERht8UF2wR+S2Ltxd55FeaXBb+D5q0zP41NZd9
1ppuZ91oOESRsnQ/zQ1a0l9Yny5de1TR5TfEqVNruU1qhjtzFcn1+LmoY5TI9nUDXK5HOyHLCG9W
X0GVOc28IWgl5pdQQqSY87ay6Ebqau0TxrCXlAV5EjY19ZPjMhkc4f5S5Wa8hHTvXEqv469zgg7m
u8JqQ9swksLlinLuCtF07Zhr+5LYwGsp4kjyLVbvGjbBaf2VWQXSDgpAO/PM1TODHq+zrqRyHYA2
Ee8xHqG70ou9kORkiZYLqlDSadgkxhnYiq0oR9716KiRQrnOjBo88/y326ckGVKifSP6wClhZMle
bjrHQsnA03qsywRYTJb3VA5OpleFqaJh/jRk+hDY4DjHTWvL6JuSUhR4EaFspYTrYF8sE3bRmvDf
fVk61e97YBQCbNJ9FzKImeesmlu2uNzNiqHHU/2BmPiddpfUHBC+4nIrdlMYCcweZ5uc08VItT7H
KHh8D8SiojjnIfisvx6FoiWBN7DK1ZXbQBpgdOmrzI8jUAgGol+HdboJ4gf3tgDGVUnJlRUqpwV0
F7ly/zPbumV22m9W/Af5LE5h5Aax+PALDavBLpFX3QH+zFc7A9PedQjg2M+aubzYGWK+uvej3piH
5YwhVEIp/wsyRYSWwr0P6QFwhjsiJGLc6IL79GNx5P4RxX1XLDQq+OI7cFQ2A1A4q/0t71PS54kq
JUMdIyLTPDRPsuLtHq0xybyq4i/L/gIHDbw0YHNA1U2ZKAvrrqEmDJ9tQmd7DCISocf9dWjdU8wr
MrdQ4MaipASgohWtU4HfDW2rbCKQsbtsfg2EsKnziDgAOSyUR2hhnH2NOgQeXoIuMoD5GR9ww70J
q5frRWHyap2nbbCxM6B4bIAHhRejYMjfuX8qNWL5Oc5HlJx7slZn3cUa3Q+XavgCScCx0S3etrHP
JrEuO+Ijaz8oSHW07B+Tf0VJgZ6ie7VT9BwoZYyilHS5qpVSCb2sr1zAZUrNKQf8i5Kx9fKahVOE
/EUvUvBdNdF9F+/C/J0oxEjrDRb774YdDoHzI39Ij6LUkGsqhjDPBKGF2accMpXxO4khnz6hjnzd
9ES+bakCt/VZNqZgywC0X3YvgwRal6WFGkBoCDriTeQGkVEv7ZL7rl1aA6QO8H0p5QIxucJyqQTC
d80zqOlL559n3QVONCqho7Evs8mbO/v0dN5SCr7pdCjQwmO9Z9MP28wR2vA+AAvqbj3j+IFQPEJB
vNGeIP2+siaueA8eMDQzA1k8lk60vpLHhz9sxvH/8+Mfb65s1lFJC+y2GWIoCB47baDd1jV85eQI
YhvjhGmGVwBWMuKVpeSm1OiQbBa+1yJZ3S2EUBnlVd6WkVkw+joKHwTZ5ViFIGWmd8pf2q+eKPbf
MmzeGgCm92ebI5vkKU4yDdZlW26nrZG5JgVY8ql+dzWV1Dgp/xVtagN5IxNiogG/iycDjF7HVkVi
Z+cvVwusQqStyhM2at/QN+aQgbePkq58osYeoeF+5M5VWJc+RcoMlQQy+d1E7ZcyblieFHVA/9v1
enTjUkNkTyRljpHOdjH/cCaSZJDhUERe6wm0iusegcbSwe0UHfaZp5z2iFCAye9mrPiEY02gyn9E
zBRWFtd6nwUaFoZolfMxS8Jk5PEFgC146oO2RAfzqknNu9hbIniyfi4lOyKbe3F9Dt8w9kwjoMIj
F2Y2v9iDfnRy8D4P38+O/EBiEl1QYr8ymQG0FHnlN2WwH4OkDIIuv3OAWgVNpJhaJ/BS1gkE3/eC
hmzq0jI0hucD7kjX6Ez+vDZje0SysRkV8qkBGv5GrZTdDiH8/PTQ+6i2AquZcwUg/YtKNKVFZv4A
W7JLSSpXafowark9aBiap3W3cHHgWg8COa8telAsIKH6fTMF7vTkhd9t77uGZxME+CCZILzIkOeA
PDIUY5xMli3dk8+t1VUufkotWCpRdqkqTJVaYuyxiF2uBT4U27C0KECiQk4IMC+G4U6h3xQN+TzE
/BDNBreH9QgFPhW7zcVwfzVIKvr7Gw+0uKTmPwOAvtXC6WuAdsEecp8r+dQw6CHdFCEbv8ZuW8gg
ejgHYywnsoacV7PehuyZUSngdpNXRmGJIVbdy2szq1WhQHKDNPhgw06MUXqWiPBEV+efo9feMZxu
MQyUIaPqp52Fr/ghBzN4Y1sCBytI2T0U+tJqGFQEFIM6hjZFYbq7ocihiv1DjFxWYvK6UVFBIlOX
Hf1pj1nDli8qZh/AlKSa1gthO7aZP8qN3tOupQRx4g1uzYLHfHzPIUrCVnFL+pdd+FjrsocYhorS
hIUoHChwpjtDRz+qyDvySO7PhYHlwb84bPQXMhEQwAVlX1dUmVc/oJOflJK+4l13cDdlwXRsocRw
qQZ+QF3w+kPBZQCYDvLV5oetLv7eSQFlu9Ot15XhCXuDB6MoS5LMGDn98Av7rQK3I8qwPx6+OtoA
bW03tNrQg+4F16+WRCHqrH09iZ4HmZZKSxMXTjM9p/fLqwFZsWgoP1wlHLgVxcANCzDI81Jnawe/
DcNUQsblgMkMA2f+RPWE/X0gyyBcCusb6EmL6ex30YPQNOXxCwz2Dln/pHOexi9faw3I22p+0Ygp
0vsnR/uyt/oLwvuFlTDPn8kRo6mjEfO8dzpfwMQwqt/j7dXeAd6OXJeD2A30XPg7DbQ7h8mJJutd
15jriTPyYK9LJUSU6InhA7xb7c2skln0oIywa7BuIMrS0vfyBbzUkE4/26Ot5tUiEiL1NTVDKvFv
Hjtcw70weJla5gRPXSOdf8OUUrRvxGJQZMs6mwGx8WQJqbHGLB8Xhp85rHyLgiBqdUEhQmSJv/xE
QZ1N94xt0NOHBs1h311hPaxP/nzEPivhvK2yd3lI+yybGUnOzfY0krOzVCVEm69rcfhwLfxomBVf
GS+WVla5vH89QIy6JTcS0Nv3GjXcOIvWlPlh74o6cK562+Xh0XbhKpDBX4almIyaSBQwnwZvpLrz
o5qqI7cftAxFo6YiH0G5Dx90h4hpug6exHCmYGnxC47G68Dt6PdTAYDY+9lYjiZHMgstQDkdwFz8
YrVnLE/jZnnAO5LCz9njnfU6ucKZ4VU4rFxT8T1mJbcvkEC04HTXbrsK2DkVauvT3denGGKeVq5c
lw+4RVleEhLmaXXi05dlgPYfgNvg1d8h0St1N/FC/kFA2+mHq3uiIFBPsXAIwY4wI0TfwpVYCk4/
MalVdgxr8JydUiLkwI56xb28/uJ4mhoWsahrWvJ7tCLagPMkK2LAyIGgk1KtQpG+JKyJiioqSyT4
IvnBd4UIJk+GdBBZu8q+h/RAbumIQJU74cu5CETJtzfa2T6ESyuOftgsFtA3Rd5HLgJonfLJm0u7
eGJvEhpEij1u5emrSUnnm/3HPQb8Xi5WpRyhKQxyRuBZR+zQ0R0Q7j0d+yyLit4zRfkLDWr7SQvw
J6EOvMTY6oKqAiJOB3ILUmGOeWOlzJg/gxCwh2YTP/IVij0Fce6c62kHBryR9DQl8xYNJ2puU8fy
KfzC7acVTv0VCSRAFecC9qyUSM4SgJIwY7aDAM0rY7y7L+2kIeDRK09Qc9t7/IPx72voIHXQQ53X
v9gNe4ly6b5FGchdSMTXLGavYQqepPgT0zsWncdajMhRMn6+lSOja4u8Sj+y/wx4XW23EMefjjFC
IGdGGBUVM4v++28pHB5RNJWhIebUH4Z1T2pB3FZZcG3YMxHEYSOauhFXpX+KLGAIh183FKjggHus
RvCXaVkH9Hs19G2PJ0XY7jm7IOpogIOv1fhjF4Asb/1n8pY/kNwHIwLOrlDVHB+bDfpqzsI8x2L+
fJqWzvaBgUurKVGvZiQ4D/6i3aHWgWzCbcBbU4z+oExM4zcvE3BrCGL7sizRNRlq8nd9qcxpHeMQ
CSkioXx66fAry4eFi12uqQegdtFTFuX9etv/nzGoCLDBRvonXeK/ClVnCWr/tK8gtHd3uaeak45E
GEgWwvSxMlAllkKZYSkKvuU52JraAmSTOgW0LXrgdCL3cCNiPq3cfbDy9QuuROS+PAbn5c6/TVES
G7nm/apKnt0Uxu8AgWv9CkyU4d5U2aCUObr0LcHExFrJKkQ6UEN4j/2+QmV81sjj04Xd1YyTCzsA
JDcmRro4kykewZ9etpHzwe+AX4u0MiktcjxUwk5rpaL/loTCCaEJ/oT1NtpRCdPWtPEKTK5mtqvs
i68EDpiFDWab5sFMo4QhdwRMq3VbHottIdlKXDdyNITrwlFCemm7dSvURPLUe+e77EyTZoxMRmyn
t+8b6sYMqSbaS4eg8y3UvR0N3vUkVv+sou8xqhA3pAIy6E5NJPNlShaAvyRBmmUcYiPrcWNlQQAF
hCDWJfY6GQQr5tVa4F188PTiKp3wzvI3wJz05Rw8s9cjzdKwAgxlTBr4tVe2/UMuqK8f0oKOWGeq
2g61450uq8D1DglZ+6jkOlI1Ps8NNblgkAwvXsQRvZkawS6gkbTpHbx+26UY4tnx5dpHxZejm0mt
W7mtMgjfGw+5c4SaVdBTNjKG23b+Unajq27yhKX0a9Je0KUarbZmKXioqAaNqR18prw85FlHpNat
7BQw1ZdtCaKP569lMpP5toeaFddD+4UqViBUnvMUzY3pBoB+NwKZ2fkfO8Zd1hTGkRP6fQo7tcMQ
dS76IqjIL8Eh+P3QIMLTPVdEjk9z/RDxoygM3zWxUJJCEZKlcnDEVl9T24j7XE1fHqV43vTeXe/u
dKT58MmCUszdE+MKY62Mr/QJDRUV7C3+uJBevtsbAwY1iblb5sX0GKzvr2BgieXRXoc0laSeG8sL
Q6vc2OLiVbGvw4jkzEJ8sOMeg3zDzd72jwJhNDLufBVswuJujXjSrzxVSAACLq3C+TcOT5I5zSMV
nQ1Q2bvuW22EW7frUdZ4LndxPaRFI2exoFHBo0hfs90/5510M70vmiMhzeqPbFJ/XXInRVt/GKtZ
NgDwWrbcK2j6PL43jEq55JZJp7ZECQcVH7/TbqbpJXNySX99P876LCbzqI3bSVwalZ9RfmpNbuts
2f33wSOOmz/ADnyebnaSahZXPPK9HAbyBDdb8VJwJUHAm2+YOcHPxOlatI4XP5XB2xXiPvNnCL6g
PJymLE7oHaH4tJ5Lx4lKD/ZRnwtfzDP+InZWQRLYU9PW6FJsZSM1KmlUj4v04TrpqpFAzMB8I3x+
TcE7AqR7RQlN8QVEW+TWpn6TFcyc3KGehWmo4z7vXGiSLQvKX5UrR2JjTVrnkgZwyAe+dVI39sNR
qacsQJSMrqKSNDh4RJEpttuVtGM1z46qnH34Ofqy7ZVmYyUPa3s4qHxaV9DIMKtuEFh9vncSkMjN
CV1YlJk9xy2k+nhemPVb++IIcl9KCXJRFdXLiz8o5aKhoD1bx4Bu9aec4CsEruSrh1yIXLc6IqPx
yw8bzT0ry1x+Dzgoo2ztXzbop5MIA5huLhoeOI0j0/A5LNELqXHUwjSC5dQi7KEExMOQt+/VbtVg
gTLrApIGbTsuGBu7DqQR/oa+gVxDl00MFxIV79B8NWRDXlh7WkojLk3AZbCvSptPlKFwQcd/rSsM
8odJxA6j6+aI1P5aSniwxqvxj9A0gluDYRHw1O0yrR0u6o92E8C6lAcZuXLwYX/3YA6oiVtKztYl
6dpu7aoyGlzbz63h7EhyRVW79jFul8voI1Ujja2NQkhq9Fea9apC7y62M+m5AqWlG1IjDzemBxdb
ub+LrX/CAVCimRCmA1lfs0uk8yYjyf5k5PQkEi1gdkfeiuHQfHEa0P4kc4vsdg1oSFFGWCtf5/SR
f9XrnSzUi9bdvknPSZk5B6jxTCx2d9p1R3ZO6ZlW9UH8vZPC2X5i5YAP9IgLCTQ7FAqngzJHxSSO
QLgjksnwxPKPDZ2ww4xsEcYPgktvpvm+MpvWsnK9pt4u6JepMYHSA3Z/Yyp0sk/F+lltbP6S/Qyp
xWPFlcg1XbvqEc//B0aT1Jtwkq5azDgaFd1m5TOCcKSWIAGeXQK+Br63Z/mhVsXjUcigs0nfzGLU
C06dBi0+tplWvAbRbbhbiLfcGBRvz85C73R16bpd9+bJ27pzvph17ezW4Qqx5smUrZ1sk69iL758
BObrhYMIYdkyp9qvbrpurVjeipHEO6VtknpJ3+PtX5wiQWtiVZOHOWQjzC1X2gV38bE0z9/25kQh
pmJJ8EkD1e+DUQde8kqQZ1yeK9re7TxPKufhp29srf5/RgJS9cwvV3fZlcPGW/A0OThg71SJa2zc
9bxqqRQj1LQZYFhnuV2bjbjckrLU253SUprmcitC3E7cux2N2nVQMovQLcr+0gzO/FBGtFZPCMj5
oFhUHnT831kH/+XUiL4+FFClE5X9zZcEMnamkQNQjeHuRPAh16lEuEssES2oP8C5v9SCxt3zyyWr
NXdx0saFCgtuaeMoa9CGVDc5o+ldQylvqxDAkR3viRzE0u8Fq2+oM/l8o40VSBX0NqLKgeMElN2U
dkIu1yztIbiucFm4Vps5gW2h9T3A9xxQbxkvnLVvo4WCtHylAXVs2p/CuXcKvGcnsLEaQ183iynV
PH93m5u4DiRe4UbnN26XBrfcLmGwQYxrtb9ofufR0138hzwxxteXL1NlJvtSglMYtSl1pKZ1k0lW
TcwIgJVbKwZCBt72kLjgcWwg+U/O7T0Kljh7gcmQmvXEkWPFCOKEN520HXYW1HLkZaikI9jWoSm0
+14je+OtSI3VaM2fQ0aEecTfIoroLlzogivENPYZA53y5HVE6Sj0uHxGJlJtJADHkNnR+MfVr/o5
vdn9HfoZN7VmtPk5EHQ/onyDD9k5NNv3XHIpVLo2kYM4xjT4oR9uQjiFhKlOCHwck1dJygbL5Z4y
G8/Ig+dSKUd+3s/mNM1VQGi8vj8rrDfW0rkcHX8aGV32tO9rstw5dM7SMCshYF54Y4n3OtnPDKgK
PkP6wKVB41+TGyHxti28iGJIwWB0fUmdtp7aAL6yLCL/nz3ZxOdWjwx094/7bTr3MYFVhQ+8KvPt
nnNpVSQy+sUmsXYfZZRHHAWZW6oRUink2/jhoHMHJtzUj5MgdR4U3COmYs4koQlUbM4N08dyIh7t
PzWkPJinS+H8q3iYPjrcI5vWJeWoh75FjkMfzWmmt2pEBrwKwihM1gF43dS7TL7SGq9s3QnDdyz9
ypX5TRLnpxNYz2nXL8W2iXLb+tmQ3yLyaBvJL4Druv3Feifhgq7/KMoX0HnqDlpGLp7wfe8CsA+a
bcd2JUgj5/Pmp1qcmlDnqtrYJ6bJ59MZso+7vxpnPCFUOJIuHnu5G83PQtpn7Wk5AkuGru+XXtdX
EMxkRZsJfTv2yD1sqnYqU3c3r301Pc9QrV/dxDekbArNfacIxxaxF+psH3NZlXdXRwAFn5+Ag3jU
suACmUDwTtZK5DH+hr9xhs7h4ek3acIxGt8XMDxI7DAx5+GVsatlcgQqiLzmNohTKcEKthaD7xmk
2HgXFzx6VUW7q1NFiidny2PHXo/vdZA1PW+S78gImuTS9w1Fhqq91lDlFP53Ex8XERlCMxClgJxn
iFIOJCI8EFS/2MsgwGyBk/ZvacYEjMGptiSXgGjgMEndeSGnInHYf1VAGEImd4lJE2GEChrQexZ2
gdPDZmX1GTQpOAav/MFlGlNyFbTpCsYVHMHUTOVwnTp2
`pragma protect end_protected
